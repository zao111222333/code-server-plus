*Version : v0p1
* .SUBCKT NHVT11LL_CKT DRN GATE SRC BULK
* +
* .ENDS
* .SUBCKT PHVT11LL_CKT DRN GATE SRC BULK
* +
* .ENDS
.SUBCKT AC1CINV2_12TH40 A B CIN CO VDD VSS
XX21 CINN XOR CO VPW NHVT11LL_CKT W=410.00n L=40.00n
XX22 BNN XNOR CO VPW NHVT11LL_CKT W=410.00n L=40.00n
XX18 CINN CIN VSS VPW NHVT11LL_CKT W=410.00n L=40.00n
XX16 BNN BN VSS VPW NHVT11LL_CKT W=410.00n L=40.00n
XX15 BN B VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX11 AN BN XNOR VPW NHVT11LL_CKT W=290.00n L=40.00n
XX12 ANN B XNOR VPW NHVT11LL_CKT W=290.00n L=40.00n
XX7 AN B XOR VPW NHVT11LL_CKT W=290.00n L=40.00n
XX5 ANN BN XOR VPW NHVT11LL_CKT W=290.00n L=40.00n
XX2 AN A VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX0 ANN AN VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX19 CINN XNOR CO VNW PHVT11LL_CKT W=500.00n L=40.00n
XX20 BNN XOR CO VNW PHVT11LL_CKT W=500.00n L=40.00n
XX17 CINN CIN VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
XX14 BNN BN VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
XX13 BN B VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX9 AN B XNOR VNW PHVT11LL_CKT W=350.00n L=40.00n
XX10 ANN BN XNOR VNW PHVT11LL_CKT W=350.00n L=40.00n
XX6 AN BN XOR VNW PHVT11LL_CKT W=350.00n L=40.00n
XX4 ANN B XOR VNW PHVT11LL_CKT W=350.00n L=40.00n
XX1 AN A VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX3 ANN AN VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS AC1CINV2_12TH40
.SUBCKT AC1CINV3_12TH40 A B CIN CO VDD VSS
XX21 CINN XOR CO VPW NHVT11LL_CKT W=0.57u L=40.00n
XX22 BNN XNOR CO VPW NHVT11LL_CKT W=0.57u L=40.00n
XX18 CINN CIN VSS VPW NHVT11LL_CKT W=0.57u L=40.00n
XX16 BNN BN VSS VPW NHVT11LL_CKT W=0.57u L=40.00n
XX15 BN B VSS VPW NHVT11LL_CKT W=0.92u L=40.00n
XX11 AN BN XNOR VPW NHVT11LL_CKT W=0.37u L=40.00n
XX12 ANN B XNOR VPW NHVT11LL_CKT W=0.37u L=40.00n
XX7 AN B XOR VPW NHVT11LL_CKT W=0.37u L=40.00n
XX5 ANN BN XOR VPW NHVT11LL_CKT W=0.37u L=40.00n
XX2 AN A VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX0 ANN AN VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX19 CINN XNOR CO VNW PHVT11LL_CKT W=0.7u L=40.00n
XX20 BNN XOR CO VNW PHVT11LL_CKT W=0.7u L=40.00n
XX17 CINN CIN VDD VNW PHVT11LL_CKT W=0.7u L=40.00n
XX14 BNN BN VDD VNW PHVT11LL_CKT W=0.7u L=40.00n
XX13 BN B VDD VNW PHVT11LL_CKT W=1.05u L=40.00n
XX9 AN B XNOR VNW PHVT11LL_CKT W=0.45u L=40.00n
XX10 ANN BN XNOR VNW PHVT11LL_CKT W=0.45u L=40.00n
XX6 AN BN XOR VNW PHVT11LL_CKT W=0.45u L=40.00n
XX4 ANN B XOR VNW PHVT11LL_CKT W=0.45u L=40.00n
XX1 AN A VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX3 ANN AN VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS AC1CINV3_12TH40
.SUBCKT AC1CINV4_12TH40 A B CIN CO VDD VSS
XX21 CINN XOR CO VPW NHVT11LL_CKT W=0.82u L=40.00n
XX22 BNN XNOR CO VPW NHVT11LL_CKT W=0.82u L=40.00n
XX18 CINN CIN VSS VPW NHVT11LL_CKT W=0.82u L=40.00n
XX16 BNN BN VSS VPW NHVT11LL_CKT W=0.82u L=40.00n
XX15 BN B VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX11 AN BN XNOR VPW NHVT11LL_CKT W=0.41u L=40.00n
XX12 ANN B XNOR VPW NHVT11LL_CKT W=0.41u L=40.00n
XX7 AN B XOR VPW NHVT11LL_CKT W=0.41u L=40.00n
XX5 ANN BN XOR VPW NHVT11LL_CKT W=0.41u L=40.00n
XX2 AN A VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX0 ANN AN VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX19 CINN XNOR CO VNW PHVT11LL_CKT W=1u L=40.00n
XX20 BNN XOR CO VNW PHVT11LL_CKT W=1u L=40.00n
XX17 CINN CIN VDD VNW PHVT11LL_CKT W=1u L=40.00n
XX14 BNN BN VDD VNW PHVT11LL_CKT W=1u L=40.00n
XX13 BN B VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX9 AN B XNOR VNW PHVT11LL_CKT W=0.5u L=40.00n
XX10 ANN BN XNOR VNW PHVT11LL_CKT W=0.5u L=40.00n
XX6 AN BN XOR VNW PHVT11LL_CKT W=0.5u L=40.00n
XX4 ANN B XOR VNW PHVT11LL_CKT W=0.5u L=40.00n
XX1 AN A VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX3 ANN AN VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS AC1CINV4_12TH40
.SUBCKT AC1CONV2_12TH40 A B CI CON VDD VSS
XX0 ANN AN VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX2 AN A VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX5 ANN BN XOR VPW NHVT11LL_CKT W=290.00n L=40.00n
XX7 AN B XOR VPW NHVT11LL_CKT W=290.00n L=40.00n
XX11 AN BN XNOR VPW NHVT11LL_CKT W=290.00n L=40.00n
XX12 ANN B XNOR VPW NHVT11LL_CKT W=290.00n L=40.00n
XX15 BN B VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX18 CIN CI VSS VPW NHVT11LL_CKT W=410.00n L=40.00n
XX21 CIN XOR CON VPW NHVT11LL_CKT W=410.00n L=40.00n
XX22 BN XNOR CON VPW NHVT11LL_CKT W=410.00n L=40.00n
XX3 ANN AN VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 AN A VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX4 ANN B XOR VNW PHVT11LL_CKT W=350.00n L=40.00n
XX6 AN BN XOR VNW PHVT11LL_CKT W=350.00n L=40.00n
XX9 AN B XNOR VNW PHVT11LL_CKT W=350.00n L=40.00n
XX10 ANN BN XNOR VNW PHVT11LL_CKT W=350.00n L=40.00n
XX13 BN B VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX17 CIN CI VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
XX19 CIN XNOR CON VNW PHVT11LL_CKT W=500.00n L=40.00n
XX20 BN XOR CON VNW PHVT11LL_CKT W=500.00n L=40.00n
.ENDS AC1CONV2_12TH40
.SUBCKT AC1CONV3_12TH40 A B CI CON VDD VSS
XX0 ANN AN VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX2 AN A VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX5 ANN BN XOR VPW NHVT11LL_CKT W=0.37u L=40.00n
XX7 AN B XOR VPW NHVT11LL_CKT W=0.37u L=40.00n
XX11 AN BN XNOR VPW NHVT11LL_CKT W=0.37u L=40.00n
XX12 ANN B XNOR VPW NHVT11LL_CKT W=0.37u L=40.00n
XX15 BN B VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX18 CIN CI VSS VPW NHVT11LL_CKT W=0.57u L=40.00n
XX21 CIN XOR CON VPW NHVT11LL_CKT W=0.57u L=40.00n
XX22 BN XNOR CON VPW NHVT11LL_CKT W=0.57u L=40.00n
XX3 ANN AN VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 AN A VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX4 ANN B XOR VNW PHVT11LL_CKT W=0.45u L=40.00n
XX6 AN BN XOR VNW PHVT11LL_CKT W=0.45u L=40.00n
XX9 AN B XNOR VNW PHVT11LL_CKT W=0.45u L=40.00n
XX10 ANN BN XNOR VNW PHVT11LL_CKT W=0.45u L=40.00n
XX13 BN B VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX17 CIN CI VDD VNW PHVT11LL_CKT W=0.7u L=40.00n
XX19 CIN XNOR CON VNW PHVT11LL_CKT W=0.7u L=40.00n
XX20 BN XOR CON VNW PHVT11LL_CKT W=0.7u L=40.00n
.ENDS AC1CONV3_12TH40
.SUBCKT AC1CONV4_12TH40 A B CI CON VDD VSS
XX0 ANN AN VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX2 AN A VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX5 ANN BN XOR VPW NHVT11LL_CKT W=0.41u L=40.00n
XX7 AN B XOR VPW NHVT11LL_CKT W=0.41u L=40.00n
XX11 AN BN XNOR VPW NHVT11LL_CKT W=0.41u L=40.00n
XX12 ANN B XNOR VPW NHVT11LL_CKT W=0.41u L=40.00n
XX15 BN B VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX18 CIN CI VSS VPW NHVT11LL_CKT W=0.82u L=40.00n
XX21 CIN XOR CON VPW NHVT11LL_CKT W=0.82u L=40.00n
XX22 BN XNOR CON VPW NHVT11LL_CKT W=0.82u L=40.00n
XX3 ANN AN VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 AN A VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX4 ANN B XOR VNW PHVT11LL_CKT W=0.5u L=40.00n
XX6 AN BN XOR VNW PHVT11LL_CKT W=0.5u L=40.00n
XX9 AN B XNOR VNW PHVT11LL_CKT W=0.5u L=40.00n
XX10 ANN BN XNOR VNW PHVT11LL_CKT W=0.5u L=40.00n
XX13 BN B VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX17 CIN CI VDD VNW PHVT11LL_CKT W=1u L=40.00n
XX19 CIN XNOR CON VNW PHVT11LL_CKT W=1u L=40.00n
XX20 BN XOR CON VNW PHVT11LL_CKT W=1u L=40.00n
.ENDS AC1CONV4_12TH40
.SUBCKT AC2CINV2_12TH40 A B CI0N CI1N CO0 CO1 VDD VSS
XX11 CO1 net62 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX10 norab ci1nn net62 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX9 nandab CI1N net62 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX8 norab ci0nn net70 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX7 nandab CI0N net70 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX6 CO0 net70 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX5 norab B VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX4 norab A VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX3 ci1nn CI1N VSS VPW NHVT11LL_CKT W=210.00n L=40.00n
XX2 net91 B VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX1 nandab A net91 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX0 ci0nn CI0N VSS VPW NHVT11LL_CKT W=210.00n L=40.00n
XX23 norab CI1N net62 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX22 nandab ci1nn net62 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX21 norab CI0N net70 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX20 nandab ci0nn net70 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX19 CO0 net70 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX18 CO1 net62 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX17 norab A net34 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX16 net34 B VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX15 nandab B VDD VNW PHVT11LL_CKT W=390.00n L=40.00n
XX14 nandab A VDD VNW PHVT11LL_CKT W=390.00n L=40.00n
XX13 ci1nn CI1N VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
XX12 ci0nn CI0N VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
.ENDS AC2CINV2_12TH40
.SUBCKT AC2CINV3_12TH40 A B CI0N CI1N CO0 CO1 VDD VSS
XX11 CO1 net62 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX10 norab ci1nn net62 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX9 nandab CI1N net62 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX8 norab ci0nn net70 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX7 nandab CI0N net70 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX6 CO0 net70 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX5 norab B VSS VPW NHVT11LL_CKT W=450.00n L=40.00n
XX4 norab A VSS VPW NHVT11LL_CKT W=450.00n L=40.00n
XX3 ci1nn CI1N VSS VPW NHVT11LL_CKT W=230.00n L=40.00n
XX2 net91 B VSS VPW NHVT11LL_CKT W=860.00n L=40.00n
XX1 nandab A net91 VPW NHVT11LL_CKT W=860.00n L=40.00n
XX0 ci0nn CI0N VSS VPW NHVT11LL_CKT W=230.00n L=40.00n
XX23 norab CI1N net62 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX22 nandab ci1nn net62 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX21 norab CI0N net70 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX20 nandab ci0nn net70 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX19 CO0 net70 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX18 CO1 net62 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX17 norab A net34 VNW PHVT11LL_CKT W=860.00n L=40.00n
XX16 net34 B VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX15 nandab B VDD VNW PHVT11LL_CKT W=550.00n L=40.00n
XX14 nandab A VDD VNW PHVT11LL_CKT W=550.00n L=40.00n
XX13 ci1nn CI1N VDD VNW PHVT11LL_CKT W=280.00n L=40.00n
XX12 ci0nn CI0N VDD VNW PHVT11LL_CKT W=280.00n L=40.00n
.ENDS AC2CINV3_12TH40
.SUBCKT AC2CINV4_12TH40 A B CI0N CI1N CO0 CO1 VDD VSS
XX11 CO1 net62 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX10 norab ci1nn net62 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX9 nandab CI1N net62 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX8 norab ci0nn net70 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX7 nandab CI0N net70 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX6 CO0 net70 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX5 norab B VSS VPW NHVT11LL_CKT W=640.00n L=40.00n
XX4 norab A VSS VPW NHVT11LL_CKT W=640.00n L=40.00n
XX3 ci1nn CI1N VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX2 net91 B VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX1 nandab A net91 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX0 ci0nn CI0N VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX23 norab CI1N net62 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX22 nandab ci1nn net62 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX21 norab CI0N net70 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX20 nandab ci0nn net70 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX19 CO0 net70 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX18 CO1 net62 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX17 norab A net34 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX16 net34 B VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX15 nandab B VDD VNW PHVT11LL_CKT W=780.00n L=40.00n
XX14 nandab A VDD VNW PHVT11LL_CKT W=780.00n L=40.00n
XX13 ci1nn CI1N VDD VNW PHVT11LL_CKT W=330.00n L=40.00n
XX12 ci0nn CI0N VDD VNW PHVT11LL_CKT W=330.00n L=40.00n
.ENDS AC2CINV4_12TH40
.SUBCKT AC2CONV2_12TH40 A B CI0 CI1 CO0N CO1N VDD VSS
XX27 orab CI1 net10 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX26 andab ci1n net10 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX25 orab CI0 net18 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX24 andab ci0n net18 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX23 CO1N net10 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX22 CO0N net18 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX21 orab norab VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX20 andab nandab VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX19 norab B VSS VPW NHVT11LL_CKT W=205.00n L=40.00n
XX18 norab A VSS VPW NHVT11LL_CKT W=205.00n L=40.00n
XX17 net47 B VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX16 nandab A net47 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX15 ci1n CI1 VSS VPW NHVT11LL_CKT W=210.00n L=40.00n
XX14 ci0n CI0 VSS VPW NHVT11LL_CKT W=210.00n L=40.00n
XX13 orab ci1n net10 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX12 andab CI1 net10 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX11 orab ci0n net18 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX10 andab CI0 net18 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX9 CO1N net10 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX8 CO0N net18 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX7 orab norab VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX6 andab nandab VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX5 norab A net98 VNW PHVT11LL_CKT W=435.00n L=40.00n
XX4 net98 B VDD VNW PHVT11LL_CKT W=435.00n L=40.00n
XX3 nandab B VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX2 nandab A VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX1 ci1n CI1 VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
XX0 ci0n CI0 VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
.ENDS AC2CONV2_12TH40
.SUBCKT AC2CONV3_12TH40 A B CI0 CI1 CO0N CO1N VDD VSS
XX27 orab CI1 net10 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX26 andab ci1n net10 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX25 orab CI0 net18 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX24 andab ci0n net18 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX23 CO1N net10 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX22 CO0N net18 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX21 orab norab VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX20 andab nandab VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX19 norab B VSS VPW NHVT11LL_CKT W=275.00n L=40.00n
XX18 norab A VSS VPW NHVT11LL_CKT W=275.00n L=40.00n
XX17 net47 B VSS VPW NHVT11LL_CKT W=450.00n L=40.00n
XX16 nandab A net47 VPW NHVT11LL_CKT W=450.00n L=40.00n
XX15 ci1n CI1 VSS VPW NHVT11LL_CKT W=230.00n L=40.00n
XX14 ci0n CI0 VSS VPW NHVT11LL_CKT W=230.00n L=40.00n
XX13 orab ci1n net10 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX12 andab CI1 net10 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX11 orab ci0n net18 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX10 andab CI0 net18 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX9 CO1N net10 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX8 CO0N net18 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX7 orab norab VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX6 andab nandab VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX5 norab A net98 VNW PHVT11LL_CKT W=580.00n L=40.00n
XX4 net98 B VDD VNW PHVT11LL_CKT W=580.00n L=40.00n
XX3 nandab B VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX2 nandab A VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX1 ci1n CI1 VDD VNW PHVT11LL_CKT W=280.00n L=40.00n
XX0 ci0n CI0 VDD VNW PHVT11LL_CKT W=280.00n L=40.00n
.ENDS AC2CONV3_12TH40
.SUBCKT AC2CONV4_12TH40 A B CI0 CI1 CO0N CO1N VDD VSS
XX27 orab CI1 net10 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX26 andab ci1n net10 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX25 orab CI0 net18 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX24 andab ci0n net18 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX23 CO1N net10 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX22 CO0N net18 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX21 orab norab VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX20 andab nandab VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX19 norab B VSS VPW NHVT11LL_CKT W=400.0n L=40.00n
XX18 norab A VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX17 net47 B VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX16 nandab A net47 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX15 ci1n CI1 VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX14 ci0n CI0 VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX13 orab ci1n net10 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX12 andab CI1 net10 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX11 orab ci0n net18 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX10 andab CI0 net18 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX9 CO1N net10 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX8 CO0N net18 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX7 orab norab VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX6 andab nandab VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX5 norab A net98 VNW PHVT11LL_CKT W=840.00n L=40.00n
XX4 net98 B VDD VNW PHVT11LL_CKT W=840.00n L=40.00n
XX3 nandab B VDD VNW PHVT11LL_CKT W=550.00n L=40.00n
XX2 nandab A VDD VNW PHVT11LL_CKT W=550.00n L=40.00n
XX1 ci1n CI1 VDD VNW PHVT11LL_CKT W=330.00n L=40.00n
XX0 ci0n CI0 VDD VNW PHVT11LL_CKT W=330.00n L=40.00n
.ENDS AC2CONV4_12TH40
.SUBCKT ACH2CONV2_12TH40 A B CO0N CO1N VDD VSS
XX3 net21 B VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX2 CO0N A net21 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX1 CO1N B VSS VPW NHVT11LL_CKT W=290.00n L=40.00n
XX0 CO1N A VSS VPW NHVT11LL_CKT W=290.00n L=40.00n
XX7 CO1N A net8 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX6 net8 B VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX5 CO0N B VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX4 CO0N A VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
.ENDS ACH2CONV2_12TH40
.SUBCKT ACH2CONV3_12TH40 A B CO0N CO1N VDD VSS
XX3 net21 B VSS VPW NHVT11LL_CKT W=860.00n L=40.00n
XX2 CO0N A net21 VPW NHVT11LL_CKT W=860.00n L=40.00n
XX1 CO1N B VSS VPW NHVT11LL_CKT W=410.00n L=40.00n
XX0 CO1N A VSS VPW NHVT11LL_CKT W=410.00n L=40.00n
XX7 CO1N A net8 VNW PHVT11LL_CKT W=860.00n L=40.00n
XX6 net8 B VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX5 CO0N B VDD VNW PHVT11LL_CKT W=560.00n L=40.00n
XX4 CO0N A VDD VNW PHVT11LL_CKT W=560.00n L=40.00n
.ENDS ACH2CONV3_12TH40
.SUBCKT ACH2CONV4_12TH40 A B CO0N CO1N VDD VSS
XX3 net21 B VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX2 CO0N A net21 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX1 CO1N B VSS VPW NHVT11LL_CKT W=580.00n L=40.00n
XX0 CO1N A VSS VPW NHVT11LL_CKT W=580.00n L=40.00n
XX7 CO1N A net8 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX6 net8 B VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX5 CO0N B VDD VNW PHVT11LL_CKT W=800.00n L=40.00n
XX4 CO0N A VDD VNW PHVT11LL_CKT W=800.00n L=40.00n
.ENDS ACH2CONV4_12TH40
.SUBCKT AD142V2_12TH40 A B C CI CO D ICO S VDD VSS
XX16 BN B VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX78 DN D VSS VPW NHVT11LL_CKT W=310.00n L=40.00n
XX79 DNN DN VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX58 BNN BN VSS VPW NHVT11LL_CKT W=300.00n L=40.00n
XX80 DN CN CD VPW NHVT11LL_CKT W=250.00n L=40.00n
XX81 DNN C CD VPW NHVT11LL_CKT W=250.00n L=40.00n
XX86 CDN CD VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX88 net0116 CDN VSS VPW NHVT11LL_CKT W=300.00n L=40.00n
XX90 net0116 AB ABCD VPW NHVT11LL_CKT W=300.00n L=40.00n
XX91 CDN ABN ABCD VPW NHVT11LL_CKT W=300.00n L=40.00n
XX94 net0104 CI VSS VPW NHVT11LL_CKT W=330.00n L=40.00n
XX95 A2DICI ABCDN net0104 VPW NHVT11LL_CKT W=330.00n L=40.00n
XX98 ICIN CI VSS VPW NHVT11LL_CKT W=240.00n L=40.00n
XX100 ABCDN ABCD VSS VPW NHVT11LL_CKT W=440.00n L=40.00n
XX101 ABCDNN ABCDN VSS VPW NHVT11LL_CKT W=300.00n L=40.00n
XX102 ABCDN CI net083 VPW NHVT11LL_CKT W=300.00n L=40.00n
XX103 ABCDNN ICIN net083 VPW NHVT11LL_CKT W=300.00n L=40.00n
XX108 S net083 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX74 CO A2DICI net076 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX75 net076 net0152 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX66 ABN AB VSS VPW NHVT11LL_CKT W=240.00n L=40.00n
XX68 CN C VSS VPW NHVT11LL_CKT W=210.00n L=40.00n
XX64 AN A VSS VPW NHVT11LL_CKT W=240.00n L=40.00n
XX61 BN AN AB VPW NHVT11LL_CKT W=300.00n L=40.00n
XX72 net088 D VSS VPW NHVT11LL_CKT W=330.00n L=40.00n
XX73 net0152 ABCD net088 VPW NHVT11LL_CKT W=330.00n L=40.00n
XX62 BNN A AB VPW NHVT11LL_CKT W=300.00n L=40.00n
XX9 net5 C VSS VPW NHVT11LL_CKT W=300.00n L=40.00n
XX8 ICON B net5 VPW NHVT11LL_CKT W=300.00n L=40.00n
XX5 net17 B VSS VPW NHVT11LL_CKT W=300.00n L=40.00n
XX2 net17 C VSS VPW NHVT11LL_CKT W=300.00n L=40.00n
XX4 ICON A net17 VPW NHVT11LL_CKT W=300.00n L=40.00n
XX11 ICO ICON VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX26 BN B VDD VNW PHVT11LL_CKT W=460.00n L=40.00n
XX59 BNN BN VDD VNW PHVT11LL_CKT W=370.00n L=40.00n
XX82 DN D VDD VNW PHVT11LL_CKT W=380.00n L=40.00n
XX83 DNN DN VDD VNW PHVT11LL_CKT W=300.00n L=40.00n
XX84 DN C CD VNW PHVT11LL_CKT W=300.00n L=40.00n
XX85 DNN CN CD VNW PHVT11LL_CKT W=300.00n L=40.00n
XX87 CDN CD VDD VNW PHVT11LL_CKT W=460.00n L=40.00n
XX89 net0116 CDN VDD VNW PHVT11LL_CKT W=370.00n L=40.00n
XX92 net0116 ABN ABCD VNW PHVT11LL_CKT W=370.00n L=40.00n
XX93 CDN AB ABCD VNW PHVT11LL_CKT W=370.00n L=40.00n
XX96 A2DICI CI VDD VNW PHVT11LL_CKT W=210.00n L=40.00n
XX97 A2DICI ABCDN VDD VNW PHVT11LL_CKT W=210.00n L=40.00n
XX99 ICIN CI VDD VNW PHVT11LL_CKT W=270.00n L=40.00n
XX104 ABCDN ABCD VDD VNW PHVT11LL_CKT W=530.00n L=40.00n
XX105 ABCDNN ABCDN VDD VNW PHVT11LL_CKT W=370.00n L=40.00n
XX106 ABCDN ICIN net083 VNW PHVT11LL_CKT W=370.00n L=40.00n
XX107 ABCDNN CI net083 VNW PHVT11LL_CKT W=370.00n L=40.00n
XX109 S net083 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX77 CO A2DICI VDD VNW PHVT11LL_CKT W=395.00n L=40.00n
XX60 BN A AB VNW PHVT11LL_CKT W=370.00n L=40.00n
XX67 ABN AB VDD VNW PHVT11LL_CKT W=270.00n L=40.00n
XX69 CN C VDD VNW PHVT11LL_CKT W=240.00n L=40.00n
XX70 net0152 D VDD VNW PHVT11LL_CKT W=210.00n L=40.00n
XX71 net0152 ABCD VDD VNW PHVT11LL_CKT W=210.00n L=40.00n
XX63 BNN AN AB VNW PHVT11LL_CKT W=370.00n L=40.00n
XX65 AN A VDD VNW PHVT11LL_CKT W=270.00n L=40.00n
XX76 CO net0152 VDD VNW PHVT11LL_CKT W=395.00n L=40.00n
XX7 ICON B net32 VNW PHVT11LL_CKT W=360.00n L=40.00n
XX6 net32 C VDD VNW PHVT11LL_CKT W=360.00n L=40.00n
XX3 ICON A net45 VNW PHVT11LL_CKT W=360.00n L=40.00n
XX0 net45 B VDD VNW PHVT11LL_CKT W=360.00n L=40.00n
XX1 net45 C VDD VNW PHVT11LL_CKT W=360.00n L=40.00n
XX10 ICO ICON VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS AD142V2_12TH40
.SUBCKT AD142V3_12TH40 A B C CI CO D ICO S VDD VSS
XX16 BN B VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX78 DN D VSS VPW NHVT11LL_CKT W=0.37u L=40.00n
XX79 DNN DN VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX58 BNN BN VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX80 DN CN CD VPW NHVT11LL_CKT W=0.3u L=40.00n
XX81 DNN C CD VPW NHVT11LL_CKT W=0.3u L=40.00n
XX86 CDN CD VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX88 net0116 CDN VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX90 net0116 AB ABCD VPW NHVT11LL_CKT W=0.4u L=40.00n
XX91 CDN ABN ABCD VPW NHVT11LL_CKT W=0.4u L=40.00n
XX94 net0104 CI VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX95 A2DICI ABCDN net0104 VPW NHVT11LL_CKT W=0.5u L=40.00n
XX98 ICIN CI VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX100 ABCDN ABCD VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX101 ABCDNN ABCDN VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX102 ABCDN CI net083 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX103 ABCDNN ICIN net083 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX108 S net083 VSS VPW NHVT11LL_CKT W=0.76u L=40.00n
XX74 CO A2DICI net076 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX75 net076 net0152 VSS VPW NHVT11LL_CKT W=0.86u L=40.00n
XX66 ABN AB VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX68 CN C VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX64 AN A VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX61 BN AN AB VPW NHVT11LL_CKT W=0.4u L=40.00n
XX72 net088 D VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX73 net0152 ABCD net088 VPW NHVT11LL_CKT W=0.5u L=40.00n
XX62 BNN A AB VPW NHVT11LL_CKT W=0.4u L=40.00n
XX9 net5 C VSS VPW NHVT11LL_CKT W=0.375u L=40.00n
XX8 ICON B net5 VPW NHVT11LL_CKT W=0.375u L=40.00n
XX5 net17 B VSS VPW NHVT11LL_CKT W=0.375u L=40.00n
XX2 net17 C VSS VPW NHVT11LL_CKT W=0.375u L=40.00n
XX4 ICON A net17 VPW NHVT11LL_CKT W=0.375u L=40.00n
XX11 ICO ICON VSS VPW NHVT11LL_CKT W=0.76u L=40.00n
XX26 BN B VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX59 BNN BN VDD VNW PHVT11LL_CKT W=0.48u L=40.00n
XX82 DN D VDD VNW PHVT11LL_CKT W=0.45u L=40.00n
XX83 DNN DN VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX84 DN C CD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX85 DNN CN CD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX87 CDN CD VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX89 net0116 CDN VDD VNW PHVT11LL_CKT W=0.48u L=40.00n
XX92 net0116 ABN ABCD VNW PHVT11LL_CKT W=0.48u L=40.00n
XX93 CDN AB ABCD VNW PHVT11LL_CKT W=0.48u L=40.00n
XX96 A2DICI CI VDD VNW PHVT11LL_CKT W=0.32u L=40.00n
XX97 A2DICI ABCDN VDD VNW PHVT11LL_CKT W=0.32u L=40.00n
XX99 ICIN CI VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX104 ABCDN ABCD VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX105 ABCDNN ABCDN VDD VNW PHVT11LL_CKT W=0.48u L=40.00n
XX106 ABCDN ICIN net083 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX107 ABCDNN CI net083 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX109 S net083 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX77 CO A2DICI VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX60 BN A AB VNW PHVT11LL_CKT W=0.48u L=40.00n
XX67 ABN AB VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX69 CN C VDD VNW PHVT11LL_CKT W=0.27u L=40.00n
XX70 net0152 D VDD VNW PHVT11LL_CKT W=0.32u L=40.00n
XX71 net0152 ABCD VDD VNW PHVT11LL_CKT W=0.32u L=40.00n
XX63 BNN AN AB VNW PHVT11LL_CKT W=0.48u L=40.00n
XX65 AN A VDD VNW PHVT11LL_CKT W=0.325u L=40.00n
XX76 CO net0152 VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX7 ICON B net32 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX6 net32 C VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
XX3 ICON A net45 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX0 net45 B VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
XX1 net45 C VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
XX10 ICO ICON VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
.ENDS AD142V3_12TH40
.SUBCKT AD142V4_12TH40 A B C CI CO D ICO S VDD VSS
XX16 BN B VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX78 DN D VSS VPW NHVT11LL_CKT W=0.37u L=40.00n
XX79 DNN DN VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX58 BNN BN VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX80 DN CN CD VPW NHVT11LL_CKT W=0.3u L=40.00n
XX81 DNN C CD VPW NHVT11LL_CKT W=0.3u L=40.00n
XX86 CDN CD VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX88 net0116 CDN VSS VPW NHVT11LL_CKT W=0.41u L=40.00n
XX90 net0116 AB ABCD VPW NHVT11LL_CKT W=0.41u L=40.00n
XX91 CDN ABN ABCD VPW NHVT11LL_CKT W=0.41u L=40.00n
XX94 net0104 CI VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX95 A2DICI ABCDN net0104 VPW NHVT11LL_CKT W=0.61u L=40.00n
XX98 ICIN CI VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX100 ABCDN ABCD VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX101 ABCDNN ABCDN VSS VPW NHVT11LL_CKT W=0.41u L=40.00n
XX102 ABCDN CI net083 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX103 ABCDNN ICIN net083 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX108 S net083 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX74 CO A2DICI net076 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX75 net076 net0152 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX66 ABN AB VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX68 CN C VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX64 AN A VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX61 BN AN AB VPW NHVT11LL_CKT W=0.4u L=40.00n
XX72 net088 D VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX73 net0152 ABCD net088 VPW NHVT11LL_CKT W=0.61u L=40.00n
XX62 BNN A AB VPW NHVT11LL_CKT W=0.4u L=40.00n
XX9 net5 C VSS VPW NHVT11LL_CKT W=0.505u L=40.00n
XX8 ICON B net5 VPW NHVT11LL_CKT W=0.505u L=40.00n
XX5 net17 B VSS VPW NHVT11LL_CKT W=0.505u L=40.00n
XX2 net17 C VSS VPW NHVT11LL_CKT W=0.505u L=40.00n
XX4 ICON A net17 VPW NHVT11LL_CKT W=0.505u L=40.00n
XX11 ICO ICON VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX26 BN B VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX59 BNN BN VDD VNW PHVT11LL_CKT W=0.48u L=40.00n
XX82 DN D VDD VNW PHVT11LL_CKT W=0.45u L=40.00n
XX83 DNN DN VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX84 DN C CD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX85 DNN CN CD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX87 CDN CD VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX89 net0116 CDN VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX92 net0116 ABN ABCD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX93 CDN AB ABCD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX96 A2DICI CI VDD VNW PHVT11LL_CKT W=0.395u L=40.00n
XX97 A2DICI ABCDN VDD VNW PHVT11LL_CKT W=0.395u L=40.00n
XX99 ICIN CI VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX104 ABCDN ABCD VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX105 ABCDNN ABCDN VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX106 ABCDN ICIN net083 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX107 ABCDNN CI net083 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX109 S net083 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX77 CO A2DICI VDD VNW PHVT11LL_CKT W=0.79u L=40.00n
XX60 BN A AB VNW PHVT11LL_CKT W=0.48u L=40.00n
XX67 ABN AB VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX69 CN C VDD VNW PHVT11LL_CKT W=0.27u L=40.00n
XX70 net0152 D VDD VNW PHVT11LL_CKT W=0.395u L=40.00n
XX71 net0152 ABCD VDD VNW PHVT11LL_CKT W=0.395u L=40.00n
XX63 BNN AN AB VNW PHVT11LL_CKT W=0.48u L=40.00n
XX65 AN A VDD VNW PHVT11LL_CKT W=0.325u L=40.00n
XX76 CO net0152 VDD VNW PHVT11LL_CKT W=0.79u L=40.00n
XX7 ICON B net32 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX6 net32 C VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX3 ICON A net45 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net45 B VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX1 net45 C VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX10 ICO ICON VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS AD142V4_12TH40
.SUBCKT AD1CINV2_12TH40 A B CIN CO S VDD VSS
XX27 CO net319 VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX24 S net323 VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX22 CINNN CINN VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX19 CINN XOR net323 VPW NHVT11LL_CKT W=270.00n L=40.00n
XX18 CINNN XNOR net323 VPW NHVT11LL_CKT W=270.00n L=40.00n
XX15 CINNN XOR net319 VPW NHVT11LL_CKT W=270.00n L=40.00n
XX14 BN XNOR net319 VPW NHVT11LL_CKT W=270.00n L=40.00n
XX12 CINN CIN VSS VPW NHVT11LL_CKT W=390.00n L=40.00n
XX9 AN BN XNOR VPW NHVT11LL_CKT W=340.00n L=40.00n
XX8 ANN B XNOR VPW NHVT11LL_CKT W=340.00n L=40.00n
XX5 ANN BN XOR VPW NHVT11LL_CKT W=340.00n L=40.00n
XX7 AN B XOR VPW NHVT11LL_CKT W=340.00n L=40.00n
XX2 ANN AN VSS VPW NHVT11LL_CKT W=510.00n L=40.00n
XX0 BN B VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX29 AN A VSS VPW NHVT11LL_CKT W=510.00n L=40.00n
XX26 CO net319 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX25 S net323 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX23 CINNN CINN VDD VNW PHVT11LL_CKT W=320.00n L=40.00n
XX21 CINN XNOR net323 VNW PHVT11LL_CKT W=320.00n L=40.00n
XX20 CINNN XOR net323 VNW PHVT11LL_CKT W=320.00n L=40.00n
XX17 CINNN XNOR net319 VNW PHVT11LL_CKT W=320.00n L=40.00n
XX16 BN XOR net319 VNW PHVT11LL_CKT W=320.00n L=40.00n
XX13 CINN CIN VDD VNW PHVT11LL_CKT W=470.00n L=40.00n
XX11 AN B XNOR VNW PHVT11LL_CKT W=400.00n L=40.00n
XX10 ANN BN XNOR VNW PHVT11LL_CKT W=400.00n L=40.00n
XX4 ANN B XOR VNW PHVT11LL_CKT W=400.00n L=40.00n
XX6 AN BN XOR VNW PHVT11LL_CKT W=400.00n L=40.00n
XX3 ANN AN VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 BN B VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX28 AN A VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS AD1CINV2_12TH40
.SUBCKT AD1CINV3_12TH40 A B CIN CO S VDD VSS
XX27 CO net319 VSS VPW NHVT11LL_CKT W=0.76u L=40.00n
XX24 S net323 VSS VPW NHVT11LL_CKT W=0.76u L=40.00n
XX22 CINNN CINN VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX19 CINN XOR net323 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX18 CINNN XNOR net323 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX15 CINNN XOR net319 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX14 BN XNOR net319 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX12 CINN CIN VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX9 AN BN XNOR VPW NHVT11LL_CKT W=0.41u L=40.00n
XX8 ANN B XNOR VPW NHVT11LL_CKT W=0.41u L=40.00n
XX5 ANN BN XOR VPW NHVT11LL_CKT W=0.41u L=40.00n
XX7 AN B XOR VPW NHVT11LL_CKT W=0.41u L=40.00n
XX2 ANN AN VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX0 BN B VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX29 AN A VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX26 CO net319 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX25 S net323 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX23 CINNN CINN VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
XX21 CINN XNOR net323 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX20 CINNN XOR net323 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX17 CINNN XNOR net319 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX16 BN XOR net319 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX13 CINN CIN VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX11 AN B XNOR VNW PHVT11LL_CKT W=0.5u L=40.00n
XX10 ANN BN XNOR VNW PHVT11LL_CKT W=0.5u L=40.00n
XX4 ANN B XOR VNW PHVT11LL_CKT W=0.5u L=40.00n
XX6 AN BN XOR VNW PHVT11LL_CKT W=0.5u L=40.00n
XX3 ANN AN VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 BN B VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX28 AN A VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS AD1CINV3_12TH40
.SUBCKT AD1CINV4_12TH40 A B CIN CO S VDD VSS
XX27 CO net319 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX24 S net323 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX22 CINNN CINN VSS VPW NHVT11LL_CKT W=0.41u L=40.00n
XX19 CINN XOR net323 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX18 CINNN XNOR net323 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX15 CINNN XOR net319 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX14 BN XNOR net319 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX12 CINN CIN VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX9 AN BN XNOR VPW NHVT11LL_CKT W=0.41u L=40.00n
XX8 ANN B XNOR VPW NHVT11LL_CKT W=0.41u L=40.00n
XX5 ANN BN XOR VPW NHVT11LL_CKT W=0.41u L=40.00n
XX7 AN B XOR VPW NHVT11LL_CKT W=0.41u L=40.00n
XX2 ANN AN VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX0 BN B VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX29 AN A VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX26 CO net319 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX25 S net323 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX23 CINNN CINN VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX21 CINN XNOR net323 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX20 CINNN XOR net323 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX17 CINNN XNOR net319 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX16 BN XOR net319 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX13 CINN CIN VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX11 AN B XNOR VNW PHVT11LL_CKT W=0.5u L=40.00n
XX10 ANN BN XNOR VNW PHVT11LL_CKT W=0.5u L=40.00n
XX4 ANN B XOR VNW PHVT11LL_CKT W=0.5u L=40.00n
XX6 AN BN XOR VNW PHVT11LL_CKT W=0.5u L=40.00n
XX3 ANN AN VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 BN B VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX28 AN A VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS AD1CINV4_12TH40
.SUBCKT AD1CONV2_12TH40 A B CI CON S VDD VSS
XX33 CON net13 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX32 net18 CI net13 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX31 net22 cin net13 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX30 net18 norab VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX29 net22 net78 VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX28 net26 B VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX27 net78 A net26 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX26 cin CI VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX25 S net49 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX24 xn cin net49 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX23 xo CI net49 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX22 xn xo VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX21 net54 B VSS VPW NHVT11LL_CKT W=430.00n L=40.00n
XX20 xo A net54 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX19 xo norab VSS VPW NHVT11LL_CKT W=260.00n L=40.00n
XX18 norab B VSS VPW NHVT11LL_CKT W=300.00n L=40.00n
XX16 norab A VSS VPW NHVT11LL_CKT W=300.00n L=40.00n
XX17 cin CI VDD VNW PHVT11LL_CKT W=390.00n L=40.00n
XX15 net78 A VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX14 net78 B VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX13 net22 net78 VDD VNW PHVT11LL_CKT W=390.00n L=40.00n
XX12 net18 norab VDD VNW PHVT11LL_CKT W=390.00n L=40.00n
XX11 CON net13 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX10 net18 cin net13 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX9 net22 CI net13 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX8 xo cin net49 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX7 xn CI net49 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX6 S net49 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX5 xn xo VDD VNW PHVT11LL_CKT W=390.00n L=40.00n
XX4 net129 B VDD VNW PHVT11LL_CKT W=520.00n L=40.00n
XX3 xo norab net129 VNW PHVT11LL_CKT W=520.00n L=40.00n
XX2 net129 A VDD VNW PHVT11LL_CKT W=520.00n L=40.00n
XX1 norab A net137 VNW PHVT11LL_CKT W=455.00n L=40.00n
XX0 net137 B VDD VNW PHVT11LL_CKT W=455.00n L=40.00n
.ENDS AD1CONV2_12TH40
.SUBCKT AD1CONV3_12TH40 A B CI CON S VDD VSS
XX33 CON net13 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX32 net18 CI net13 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX31 net22 cin net13 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX30 net18 norab VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX29 net22 net78 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX28 net26 B VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX27 net78 A net26 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX26 cin CI VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX25 S net49 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX24 xn cin net49 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX23 xo CI net49 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX22 xn xo VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX21 net54 B VSS VPW NHVT11LL_CKT W=460.00n L=40.00n
XX20 xo A net54 VPW NHVT11LL_CKT W=460.00n L=40.00n
XX19 xo norab VSS VPW NHVT11LL_CKT W=280.00n L=40.00n
XX18 norab B VSS VPW NHVT11LL_CKT W=325.00n L=40.00n
XX16 norab A VSS VPW NHVT11LL_CKT W=325.00n L=40.00n
XX17 cin CI VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX15 net78 A VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
XX14 net78 B VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
XX13 net22 net78 VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX12 net18 norab VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX11 CON net13 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX10 net18 cin net13 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX9 net22 CI net13 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX8 xo cin net49 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX7 xn CI net49 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX6 S net49 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX5 xn xo VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX4 net129 B VDD VNW PHVT11LL_CKT W=560.00n L=40.00n
XX3 xo norab net129 VNW PHVT11LL_CKT W=560.00n L=40.00n
XX2 net129 A VDD VNW PHVT11LL_CKT W=560.00n L=40.00n
XX1 norab A net137 VNW PHVT11LL_CKT W=495.00n L=40.00n
XX0 net137 B VDD VNW PHVT11LL_CKT W=495.00n L=40.00n
.ENDS AD1CONV3_12TH40
.SUBCKT AD1CONV4_12TH40 A B CI CON S VDD VSS
XX33 CON net13 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX32 net18 CI net13 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX31 net22 cin net13 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX30 net18 norab VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX29 net22 net78 VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX28 net26 B VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX27 net78 A net26 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX26 cin CI VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX25 S net49 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX24 xn cin net49 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX23 xo CI net49 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX22 xn xo VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX21 net54 B VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX20 xo A net54 VPW NHVT11LL_CKT W=500.00n L=40.00n
XX19 xo norab VSS VPW NHVT11LL_CKT W=300.00n L=40.00n
XX18 norab B VSS VPW NHVT11LL_CKT W=370.00n L=40.00n
XX16 norab A VSS VPW NHVT11LL_CKT W=370.00n L=40.00n
XX17 cin CI VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
XX15 net78 A VDD VNW PHVT11LL_CKT W=355.00n L=40.00n
XX14 net78 B VDD VNW PHVT11LL_CKT W=355.00n L=40.00n
XX13 net22 net78 VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
XX12 net18 norab VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
XX11 CON net13 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX10 net18 cin net13 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX9 net22 CI net13 VNW PHVT11LL_CKT W=465.00n L=40.00n
XX8 xo cin net49 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX7 xn CI net49 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX6 S net49 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX5 xn xo VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
XX4 net129 B VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX3 xo norab net129 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX2 net129 A VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 norab A net137 VNW PHVT11LL_CKT W=560.00n L=40.00n
XX0 net137 B VDD VNW PHVT11LL_CKT W=560.00n L=40.00n
.ENDS AD1CONV4_12TH40
.SUBCKT AD1V2C_12TH40 A B CI CO S VDD VSS
XX25 S net45 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX23 net0187 CI VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX22 net0187 B VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX20 net0179 B VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX19 net0183 A net0179 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX21 net0187 A VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX18 net45 CI net0183 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX17 net45 net0129 net0187 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX9 net0129 A net49 VPW NHVT11LL_CKT W=270.00n L=40.00n
XX8 net49 B VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX4 CO net0129 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX3 net0129 CI net61 VPW NHVT11LL_CKT W=270.00n L=40.00n
XX2 net61 B VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX29 net61 A VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX24 S net45 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX16 net45 CI net0118 VNW PHVT11LL_CKT W=425.00n L=40.00n
XX14 net0126 B VDD VNW PHVT11LL_CKT W=425.00n L=40.00n
XX15 net0118 A net0126 VNW PHVT11LL_CKT W=425.00n L=40.00n
XX13 net45 net0129 net9 VNW PHVT11LL_CKT W=425.00n L=40.00n
XX12 net9 CI VDD VNW PHVT11LL_CKT W=425.00n L=40.00n
XX11 net9 A VDD VNW PHVT11LL_CKT W=425.00n L=40.00n
XX10 net9 B VDD VNW PHVT11LL_CKT W=425.00n L=40.00n
XX7 net0129 A net24 VNW PHVT11LL_CKT W=325.00n L=40.00n
XX6 net24 B VDD VNW PHVT11LL_CKT W=325.00n L=40.00n
XX5 CO net0129 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 net0129 CI net37 VNW PHVT11LL_CKT W=325.00n L=40.00n
XX0 net37 B VDD VNW PHVT11LL_CKT W=325.00n L=40.00n
XX28 net37 A VDD VNW PHVT11LL_CKT W=325.00n L=40.00n
.ENDS AD1V2C_12TH40
.SUBCKT AD1V2R_12TH40 A B CI CO S VDD VSS
XX2 cin CI VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX25 S net41 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX7 xo A net54 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX23 norab CI net21 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX21 net106 cin net21 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX14 net26 B VSS VPW NHVT11LL_CKT W=450.00n L=40.00n
XX27 CO net21 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX0 norab A VSS VPW NHVT11LL_CKT W=490.00n L=40.00n
XX19 xo CI net41 VPW NHVT11LL_CKT W=320.00n L=40.00n
XXN1 xo norab VSS VPW NHVT11LL_CKT W=260.00n L=40.00n
XX11 xn xo VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX5 norab B VSS VPW NHVT11LL_CKT W=490.00n L=40.00n
XX8 net54 B VSS VPW NHVT11LL_CKT W=430.00n L=40.00n
XX13 net106 A net26 VPW NHVT11LL_CKT W=450.00n L=40.00n
XX17 xn cin net41 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX20 net106 CI net21 VNW PHVT11LL_CKT W=390.00n L=40.00n
XXP1 net81 A VDD VNW PHVT11LL_CKT W=520.00n L=40.00n
XX4 norab A net77 VNW PHVT11LL_CKT W=880.00n L=40.00n
XX6 xo norab net81 VNW PHVT11LL_CKT W=520.00n L=40.00n
XX3 net77 B VDD VNW PHVT11LL_CKT W=880.00n L=40.00n
XX24 S net41 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX9 net81 B VDD VNW PHVT11LL_CKT W=520.00n L=40.00n
XX18 xo cin net41 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX10 xn xo VDD VNW PHVT11LL_CKT W=390.00n L=40.00n
XX22 norab cin net21 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX12 net106 A VDD VNW PHVT11LL_CKT W=390.00n L=40.00n
XX26 CO net21 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX15 net106 B VDD VNW PHVT11LL_CKT W=390.00n L=40.00n
XX16 xn CI net41 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX1 cin CI VDD VNW PHVT11LL_CKT W=390.00n L=40.00n
.ENDS AD1V2R_12TH40
.SUBCKT AD1V2T_12TH40 A B CI CO S VDD VSS
XX19 xn xo VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX23 xo CI net13 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX21 xn cin net13 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX25 S net13 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX17 CO net53 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX1 cin CI VSS VPW NHVT11LL_CKT W=480.00n L=40.00n
XX14 net30 B VSS VPW NHVT11LL_CKT W=430.00n L=40.00n
XX13 xo A net30 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX4 net38 A VSS VPW NHVT11LL_CKT W=200.00n L=40.00n
XX7 net38 B VSS VPW NHVT11LL_CKT W=200.00n L=40.00n
XXN1 xo net38 VSS VPW NHVT11LL_CKT W=260.00n L=40.00n
XX11 net58 xn net53 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX9 cin xo net53 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX3 net58 B VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX8 cin xn net53 VNW PHVT11LL_CKT W=390.00n L=40.00n
XXP1 net93 A VDD VNW PHVT11LL_CKT W=520.00n L=40.00n
XX6 net38 A net73 VNW PHVT11LL_CKT W=345.00n L=40.00n
XX18 xn xo VDD VNW PHVT11LL_CKT W=390.00n L=40.00n
XX10 net58 xo net53 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX16 CO net53 VDD VNW PHVT11LL_CKT W=610n L=40.00n
XX20 xn CI net13 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX12 xo net38 net93 VNW PHVT11LL_CKT W=520.00n L=40.00n
XX5 net73 B VDD VNW PHVT11LL_CKT W=345.00n L=40.00n
XX24 S net13 VDD VNW PHVT11LL_CKT W=610n L=40.00n
XX15 net93 B VDD VNW PHVT11LL_CKT W=520.00n L=40.00n
XX22 xo cin net13 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX2 net58 B VDD VNW PHVT11LL_CKT W=390.00n L=40.00n
XX0 cin CI VDD VNW PHVT11LL_CKT W=585.00n L=40.00n
.ENDS AD1V2T_12TH40
.SUBCKT AD1V2_12TH40 A B CI CO S VDD VSS
XX27 CO net059 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX24 S net055 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX22 CINN CIN VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX19 CINN XOR net055 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX18 CIN XNOR net055 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX15 CIN XOR net059 VPW NHVT11LL_CKT W=270.00n L=40.00n
XX14 BN XNOR net059 VPW NHVT11LL_CKT W=270.00n L=40.00n
XX12 CIN CI VSS VPW NHVT11LL_CKT W=390.00n L=40.00n
XX9 AN BN XNOR VPW NHVT11LL_CKT W=340.00n L=40.00n
XX8 ANN B XNOR VPW NHVT11LL_CKT W=340.00n L=40.00n
XX5 ANN BN XOR VPW NHVT11LL_CKT W=340.00n L=40.00n
XX7 AN B XOR VPW NHVT11LL_CKT W=340.00n L=40.00n
XX2 ANN AN VSS VPW NHVT11LL_CKT W=510.00n L=40.00n
XX0 BN B VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX29 AN A VSS VPW NHVT11LL_CKT W=510.00n L=40.00n
XX26 CO net059 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX25 S net055 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX23 CINN CIN VDD VNW PHVT11LL_CKT W=320.00n L=40.00n
XX21 CINN XNOR net055 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX20 CIN XOR net055 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX17 CIN XNOR net059 VNW PHVT11LL_CKT W=320.00n L=40.00n
XX16 BN XOR net059 VNW PHVT11LL_CKT W=320.00n L=40.00n
XX13 CIN CI VDD VNW PHVT11LL_CKT W=470.00n L=40.00n
XX11 AN B XNOR VNW PHVT11LL_CKT W=400.00n L=40.00n
XX10 ANN BN XNOR VNW PHVT11LL_CKT W=400.00n L=40.00n
XX4 ANN B XOR VNW PHVT11LL_CKT W=400.00n L=40.00n
XX6 AN BN XOR VNW PHVT11LL_CKT W=400.00n L=40.00n
XX3 ANN AN VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 BN B VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX28 AN A VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS AD1V2_12TH40
.SUBCKT AD1V3C_12TH40 A B CI CO S VDD VSS
XX25 S net45 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX23 net0187 CI VSS VPW NHVT11LL_CKT W=0.41u L=40.00n
XX22 net0187 B VSS VPW NHVT11LL_CKT W=0.41u L=40.00n
XX20 net0179 B VSS VPW NHVT11LL_CKT W=0.41u L=40.00n
XX19 net0183 A net0179 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX21 net0187 A VSS VPW NHVT11LL_CKT W=0.41u L=40.00n
XX18 net45 CI net0183 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX17 net45 net0129 net0187 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX9 net0129 A net49 VPW NHVT11LL_CKT W=0.35u L=40.00n
XX8 net49 B VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX4 CO net0129 VSS VPW NHVT11LL_CKT W=0.75u L=40.00n
XX3 net0129 CI net61 VPW NHVT11LL_CKT W=0.35u L=40.00n
XX2 net61 B VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX29 net61 A VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX24 S net45 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX16 net45 CI net0118 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX14 net0126 B VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX15 net0118 A net0126 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX13 net45 net0129 net9 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX12 net9 CI VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX11 net9 A VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX10 net9 B VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX7 net0129 A net24 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX6 net24 B VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX5 CO net0129 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX1 net0129 CI net37 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX0 net37 B VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX28 net37 A VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
.ENDS AD1V3C_12TH40
.SUBCKT AD1V3R_12TH40 A B CI CO S VDD VSS
XX2 cin CI VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX25 S net41 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX7 xo A net54 VPW NHVT11LL_CKT W=460.00n L=40.00n
XX23 norab CI net21 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX21 net106 cin net21 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX14 net26 B VSS VPW NHVT11LL_CKT W=470.00n L=40.00n
XX27 CO net21 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX0 norab A VSS VPW NHVT11LL_CKT W=530.00n L=40.00n
XX19 xo CI net41 VPW NHVT11LL_CKT W=350.00n L=40.00n
XXN1 xo norab VSS VPW NHVT11LL_CKT W=280.00n L=40.00n
XX11 xn xo VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX5 norab B VSS VPW NHVT11LL_CKT W=530.00n L=40.00n
XX8 net54 B VSS VPW NHVT11LL_CKT W=460.00n L=40.00n
XX13 net106 A net26 VPW NHVT11LL_CKT W=470.00n L=40.00n
XX17 xn cin net41 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX20 net106 CI net21 VNW PHVT11LL_CKT W=420.00n L=40.00n
XXP1 net81 A VDD VNW PHVT11LL_CKT W=560.00n L=40.00n
XX4 norab A net77 VNW PHVT11LL_CKT W=950.00n L=40.00n
XX6 xo norab net81 VNW PHVT11LL_CKT W=560.00n L=40.00n
XX3 net77 B VDD VNW PHVT11LL_CKT W=950.00n L=40.00n
XX24 S net41 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX9 net81 B VDD VNW PHVT11LL_CKT W=560.00n L=40.00n
XX18 xo cin net41 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX10 xn xo VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX22 norab cin net21 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX12 net106 A VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX26 CO net21 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX15 net106 B VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX16 xn CI net41 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX1 cin CI VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
.ENDS AD1V3R_12TH40
.SUBCKT AD1V3T_12TH40 A B CI CO S VDD VSS
XX19 xn xo VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX23 xo CI net13 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX21 xn cin net13 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX25 S net13 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX17 CO net53 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX1 cin CI VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX14 net30 B VSS VPW NHVT11LL_CKT W=460.00n L=40.00n
XX13 xo A net30 VPW NHVT11LL_CKT W=460.00n L=40.00n
XX4 net38 A VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX7 net38 B VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XXN1 xo net38 VSS VPW NHVT11LL_CKT W=280.00n L=40.00n
XX11 net58 xn net53 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX9 cin xo net53 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX3 net58 B VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX8 cin xn net53 VNW PHVT11LL_CKT W=420.00n L=40.00n
XXP1 net93 A VDD VNW PHVT11LL_CKT W=560.00n L=40.00n
XX6 net38 A net73 VNW PHVT11LL_CKT W=380.00n L=40.00n
XX18 xn xo VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX10 net58 xo net53 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX16 CO net53 VDD VNW PHVT11LL_CKT W=860n L=40.00n
XX20 xn CI net13 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX12 xo net38 net93 VNW PHVT11LL_CKT W=560.00n L=40.00n
XX5 net73 B VDD VNW PHVT11LL_CKT W=380.00n L=40.00n
XX24 S net13 VDD VNW PHVT11LL_CKT W=860n L=40.00n
XX15 net93 B VDD VNW PHVT11LL_CKT W=560.00n L=40.00n
XX22 xo cin net13 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX2 net58 B VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX0 cin CI VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS AD1V3T_12TH40
.SUBCKT AD1V3_12TH40 A B CI CO S VDD VSS
XX27 CO net059 VSS VPW NHVT11LL_CKT W=0.75u L=40.00n
XX24 S net055 VSS VPW NHVT11LL_CKT W=0.75u L=40.00n
XX22 CINN CIN VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX19 CINN XOR net055 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX18 CIN XNOR net055 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX15 CIN XOR net059 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX14 BN XNOR net059 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX12 CIN CI VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX9 AN BN XNOR VPW NHVT11LL_CKT W=0.41u L=40.00n
XX8 ANN B XNOR VPW NHVT11LL_CKT W=0.41u L=40.00n
XX5 ANN BN XOR VPW NHVT11LL_CKT W=0.41u L=40.00n
XX7 AN B XOR VPW NHVT11LL_CKT W=0.41u L=40.00n
XX2 ANN AN VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX0 BN B VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX29 AN A VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX26 CO net059 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX25 S net055 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX23 CINN CIN VDD VNW PHVT11LL_CKT W=0.465u L=40.00n
XX21 CINN XNOR net055 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX20 CIN XOR net055 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX17 CIN XNOR net059 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX16 BN XOR net059 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX13 CIN CI VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX11 AN B XNOR VNW PHVT11LL_CKT W=0.5u L=40.00n
XX10 ANN BN XNOR VNW PHVT11LL_CKT W=0.5u L=40.00n
XX4 ANN B XOR VNW PHVT11LL_CKT W=0.5u L=40.00n
XX6 AN BN XOR VNW PHVT11LL_CKT W=0.5u L=40.00n
XX3 ANN AN VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 BN B VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX28 AN A VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS AD1V3_12TH40
.SUBCKT AD1V4C_12TH40 A B CI CO S VDD VSS
XX25 S net45 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX23 net0187 CI VSS VPW NHVT11LL_CKT W=0.41u L=40.00n
XX22 net0187 B VSS VPW NHVT11LL_CKT W=0.41u L=40.00n
XX20 net0179 B VSS VPW NHVT11LL_CKT W=0.41u L=40.00n
XX19 net0183 A net0179 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX21 net0187 A VSS VPW NHVT11LL_CKT W=0.41u L=40.00n
XX18 net45 CI net0183 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX17 net45 net0129 net0187 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX9 net0129 A net49 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX8 net49 B VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX4 CO net0129 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX3 net0129 CI net61 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX2 net61 B VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX29 net61 A VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX24 S net45 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX16 net45 CI net0118 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX14 net0126 B VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX15 net0118 A net0126 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX13 net45 net0129 net9 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX12 net9 CI VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX11 net9 A VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX10 net9 B VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX7 net0129 A net24 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX6 net24 B VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX5 CO net0129 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 net0129 CI net37 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX0 net37 B VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX28 net37 A VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
.ENDS AD1V4C_12TH40
.SUBCKT AD1V4R_12TH40 A B CI CO S VDD VSS
XX2 cin CI VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX25 S net41 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX7 xo A net54 VPW NHVT11LL_CKT W=500.00n L=40.00n
XX23 norab CI net21 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX21 net106 cin net21 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX14 net26 B VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX27 CO net21 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX0 norab A VSS VPW NHVT11LL_CKT W=570.00n L=40.00n
XX19 xo CI net41 VPW NHVT11LL_CKT W=400.00n L=40.00n
XXN1 xo norab VSS VPW NHVT11LL_CKT W=300.00n L=40.00n
XX11 xn xo VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX5 norab B VSS VPW NHVT11LL_CKT W=570.00n L=40.00n
XX8 net54 B VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX13 net106 A net26 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX17 xn cin net41 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX20 net106 CI net21 VNW PHVT11LL_CKT W=500.00n L=40.00n
XXP1 net81 A VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX4 norab A net77 VNW PHVT11LL_CKT W=1.03u L=40.00n
XX6 xo norab net81 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX3 net77 B VDD VNW PHVT11LL_CKT W=1.03u L=40.00n
XX24 S net41 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX9 net81 B VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX18 xo cin net41 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX10 xn xo VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
XX22 norab cin net21 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX12 net106 A VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
XX26 CO net21 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX15 net106 B VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
XX16 xn CI net41 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX1 cin CI VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
.ENDS AD1V4R_12TH40
.SUBCKT AD1V4T_12TH40 A B CI CO S VDD VSS
XX19 xn xo VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX23 xo CI net13 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX21 xn cin net13 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX25 S net13 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX17 CO net53 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX1 cin CI VSS VPW NHVT11LL_CKT W=600.00n L=40.00n
XX14 net30 B VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX13 xo A net30 VPW NHVT11LL_CKT W=500.00n L=40.00n
XX4 net38 A VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX7 net38 B VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XXN1 xo net38 VSS VPW NHVT11LL_CKT W=300.00n L=40.00n
XX11 net58 xn net53 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX9 cin xo net53 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX3 net58 B VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX8 cin xn net53 VNW PHVT11LL_CKT W=500.00n L=40.00n
XXP1 net93 A VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX6 net38 A net73 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX18 xn xo VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
XX10 net58 xo net53 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX16 CO net53 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX20 xn CI net13 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX12 xo net38 net93 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX5 net73 B VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX24 S net13 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX15 net93 B VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX22 xo cin net13 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX2 net58 B VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
XX0 cin CI VDD VNW PHVT11LL_CKT W=750.00n L=40.00n
.ENDS AD1V4T_12TH40
.SUBCKT AD1V4_12TH40 A B CI CO S VDD VSS
XX27 CO net059 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX24 S net055 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX22 CINN CIN VSS VPW NHVT11LL_CKT W=0.41u L=40.00n
XX19 CINN XOR net055 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX18 CIN XNOR net055 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX15 CIN XOR net059 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX14 BN XNOR net059 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX12 CIN CI VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX9 AN BN XNOR VPW NHVT11LL_CKT W=0.41u L=40.00n
XX8 ANN B XNOR VPW NHVT11LL_CKT W=0.41u L=40.00n
XX5 ANN BN XOR VPW NHVT11LL_CKT W=0.41u L=40.00n
XX7 AN B XOR VPW NHVT11LL_CKT W=0.41u L=40.00n
XX2 ANN AN VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX0 BN B VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX29 AN A VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX26 CO net059 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX25 S net055 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX23 CINN CIN VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX21 CINN XNOR net055 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX20 CIN XOR net055 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX17 CIN XNOR net059 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX16 BN XOR net059 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX13 CIN CI VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX11 AN B XNOR VNW PHVT11LL_CKT W=0.5u L=40.00n
XX10 ANN BN XNOR VNW PHVT11LL_CKT W=0.5u L=40.00n
XX4 ANN B XOR VNW PHVT11LL_CKT W=0.5u L=40.00n
XX6 AN BN XOR VNW PHVT11LL_CKT W=0.5u L=40.00n
XX3 ANN AN VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 BN B VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX28 AN A VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS AD1V4_12TH40
.SUBCKT AD2CSCINV2_12TH40 A B CI0N CI1N CO0 CO1 CS S VDD VSS
XX3 ci1nn CI1N VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX1 ci0nn CI0N VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX7 ci0 CI0N VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX5 csn CS VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX15 ci1 CI1N VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX29 norab ci0nn net32 VPW NHVT11LL_CKT W=0.35u L=40.00n
XX27 nandab CI0N net32 VPW NHVT11LL_CKT W=0.35u L=40.00n
XX19 net37 B VSS VPW NHVT11LL_CKT W=0.86u L=40.00n
XX18 nandab A net37 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX33 CO0 net32 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX51 CO1 net56 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX45 norab ci1nn net56 VPW NHVT11LL_CKT W=0.35u L=40.00n
XX43 nandab CI1N net56 VPW NHVT11LL_CKT W=0.35u L=40.00n
XX41 net89 CI1N net64 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX49 net64 CS net68 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX39 net93 ci1 net64 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX47 net80 csn net68 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX37 net89 CI0N net80 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX35 net93 ci0 net80 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX53 S net68 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX31 net89 net93 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX25 net93 net181 VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX23 net97 net105 VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX22 net181 nandab net97 VPW NHVT11LL_CKT W=0.32u L=40.00n
XX13 net105 norab VSS VPW NHVT11LL_CKT W=0.235u L=40.00n
XX11 norab B VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX8 norab A VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX44 norab CI1N net56 VNW PHVT11LL_CKT W=0.42u L=40.00n
XX42 nandab ci1nn net56 VNW PHVT11LL_CKT W=0.42u L=40.00n
XX50 CO1 net56 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX32 CO0 net32 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX28 norab CI0N net32 VNW PHVT11LL_CKT W=0.42u L=40.00n
XX26 nandab ci0nn net32 VNW PHVT11LL_CKT W=0.42u L=40.00n
XX20 nandab B VDD VNW PHVT11LL_CKT W=0.76u L=40.00n
XX17 nandab A VDD VNW PHVT11LL_CKT W=0.76u L=40.00n
XX14 ci1 CI1N VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX6 ci0 CI0N VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX4 csn CS VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX2 ci1nn CI1N VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX0 ci0nn CI0N VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX12 net105 norab VDD VNW PHVT11LL_CKT W=0.285u L=40.00n
XX10 norab A net176 VNW PHVT11LL_CKT W=0.86u L=40.00n
XX9 net176 B VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX16 net181 nandab VDD VNW PHVT11LL_CKT W=0.285u L=40.00n
XX21 net181 net105 VDD VNW PHVT11LL_CKT W=0.285u L=40.00n
XX24 net93 net181 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX30 net89 net93 VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX40 net89 ci1 net64 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX46 net80 CS net68 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX34 net93 CI0N net80 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX52 S net68 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX48 net64 csn net68 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX38 net93 CI1N net64 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX36 net89 ci0 net80 VNW PHVT11LL_CKT W=0.5u L=40.00n
.ENDS AD2CSCINV2_12TH40
.SUBCKT AD2CSCINV3_12TH40 A B CI0N CI1N CO0 CO1 CS S VDD VSS
XX3 ci1nn CI1N VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX1 ci0nn CI0N VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX7 ci0 CI0N VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX5 csn CS VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX15 ci1 CI1N VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX29 norab ci0nn net32 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX27 nandab CI0N net32 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX19 net37 B VSS VPW NHVT11LL_CKT W=860.00n L=40.00n
XX18 nandab A net37 VPW NHVT11LL_CKT W=860.00n L=40.00n
XX33 CO0 net32 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX51 CO1 net56 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX45 norab ci1nn net56 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX43 nandab CI1N net56 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX41 net89 CI1N net64 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX49 net64 CS net68 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX39 net93 ci1 net64 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX47 net80 csn net68 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX37 net89 CI0N net80 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX35 net93 ci0 net80 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX53 S net68 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX31 net89 net93 VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX25 net93 net181 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX23 net97 net105 VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX22 net181 nandab net97 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX13 net105 norab VSS VPW NHVT11LL_CKT W=235.00n L=40.00n
XX11 norab B VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX8 norab A VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX44 norab CI1N net56 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX42 nandab ci1nn net56 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX50 CO1 net56 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX32 CO0 net32 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX28 norab CI0N net32 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX26 nandab ci0nn net32 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX20 nandab B VDD VNW PHVT11LL_CKT W=760.00n L=40.00n
XX17 nandab A VDD VNW PHVT11LL_CKT W=760.00n L=40.00n
XX14 ci1 CI1N VDD VNW PHVT11LL_CKT W=330.00n L=40.00n
XX6 ci0 CI0N VDD VNW PHVT11LL_CKT W=330.00n L=40.00n
XX4 csn CS VDD VNW PHVT11LL_CKT W=330.00n L=40.00n
XX2 ci1nn CI1N VDD VNW PHVT11LL_CKT W=330.00n L=40.00n
XX0 ci0nn CI0N VDD VNW PHVT11LL_CKT W=330.00n L=40.00n
XX12 net105 norab VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX10 norab A net176 VNW PHVT11LL_CKT W=860.00n L=40.00n
XX9 net176 B VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX16 net181 nandab VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX21 net181 net105 VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX24 net93 net181 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX30 net89 net93 VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
XX40 net89 ci1 net64 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX46 net80 CS net68 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX34 net93 CI0N net80 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX52 S net68 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX48 net64 csn net68 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX38 net93 CI1N net64 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX36 net89 ci0 net80 VNW PHVT11LL_CKT W=500.00n L=40.00n
.ENDS AD2CSCINV3_12TH40
.SUBCKT AD2CSCINV4_12TH40 A B CI0N CI1N CO0 CO1 CS S VDD VSS
XX3 ci1nn CI1N VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX1 ci0nn CI0N VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX7 ci0 CI0N VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX5 csn CS VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX15 ci1 CI1N VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX29 norab ci0nn net32 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX27 nandab CI0N net32 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX19 net37 B VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX18 nandab A net37 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX33 CO0 net32 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX51 CO1 net56 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX45 norab ci1nn net56 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX43 nandab CI1N net56 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX41 net89 CI1N net64 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX49 net64 CS net68 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX39 net93 ci1 net64 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX47 net80 csn net68 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX37 net89 CI0N net80 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX35 net93 ci0 net80 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX53 S net68 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX31 net89 net93 VSS VPW NHVT11LL_CKT W=690.00n L=40.00n
XX25 net93 net181 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX23 net97 net105 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX22 net181 nandab net97 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX13 net105 norab VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX11 norab B VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX8 norab A VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX44 norab CI1N net56 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX42 nandab ci1nn net56 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX50 CO1 net56 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX32 CO0 net32 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX28 norab CI0N net32 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX26 nandab ci0nn net32 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX20 nandab B VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX17 nandab A VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX14 ci1 CI1N VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX6 ci0 CI0N VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX4 csn CS VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX2 ci1nn CI1N VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX0 ci0nn CI0N VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX12 net105 norab VDD VNW PHVT11LL_CKT W=330.00n L=40.00n
XX10 norab A net176 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX9 net176 B VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX16 net181 nandab VDD VNW PHVT11LL_CKT W=550.00n L=40.00n
XX21 net181 net105 VDD VNW PHVT11LL_CKT W=550.00n L=40.00n
XX24 net93 net181 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX30 net89 net93 VDD VNW PHVT11LL_CKT W=870.00n L=40.00n
XX40 net89 ci1 net64 VNW PHVT11LL_CKT W=870.00n L=40.00n
XX46 net80 CS net68 VNW PHVT11LL_CKT W=870.00n L=40.00n
XX34 net93 CI0N net80 VNW PHVT11LL_CKT W=870.00n L=40.00n
XX52 S net68 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX48 net64 csn net68 VNW PHVT11LL_CKT W=870.00n L=40.00n
XX38 net93 CI1N net64 VNW PHVT11LL_CKT W=870.00n L=40.00n
XX36 net89 ci0 net80 VNW PHVT11LL_CKT W=870.00n L=40.00n
.ENDS AD2CSCINV4_12TH40
.SUBCKT AD2CSCONV2_12TH40 A B CI0 CI1 CO0N CO1N CS S VDD VSS
XX3 ci1nnn CI1 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX1 ci0nnn CI0 VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX9 csn CS VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX7 ci1n CI1 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX5 ci0n CI0 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX17 net141 B VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX16 nandab A net141 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX31 orab CI0 net152 VPW NHVT11LL_CKT W=0.34u L=40.00n
XX29 andab ci0n net152 VPW NHVT11LL_CKT W=0.34u L=40.00n
XX25 orab norab VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX23 andab nandab VSS VPW NHVT11LL_CKT W=0.325u L=40.00n
XX35 CO0N net152 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX55 CO1N net176 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX47 orab CI1 net176 VPW NHVT11LL_CKT W=0.325u L=40.00n
XX45 andab ci1n net176 VPW NHVT11LL_CKT W=0.325u L=40.00n
XX43 net213 CI1 net184 VPW NHVT11LL_CKT W=0.265u L=40.00n
XX51 net184 CS net188 VPW NHVT11LL_CKT W=0.325u L=40.00n
XX41 net209 ci1nnn net184 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX49 net200 csn net188 VPW NHVT11LL_CKT W=0.325u L=40.00n
XX39 net213 CI0 net200 VPW NHVT11LL_CKT W=0.21u L=40.00n
XX37 net209 ci0nnn net200 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX53 S net188 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX33 net209 net213 VSS VPW NHVT11LL_CKT W=340.00n L=40.00n
XX27 net213 net37 VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX21 net217 orab VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX20 net37 nandab net217 VPW NHVT11LL_CKT W=0.34u L=40.00n
XX13 norab B VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX10 norab A VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX42 net213 ci1nnn net184 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX40 net209 CI1 net184 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX38 net213 ci0nnn net200 VNW PHVT11LL_CKT W=0.41u L=40.00n
XX36 net209 CI0 net200 VNW PHVT11LL_CKT W=0.41u L=40.00n
XX32 net209 net213 VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX26 net213 net37 VDD VNW PHVT11LL_CKT W=0.41u L=40.00n
XX19 net37 orab VDD VNW PHVT11LL_CKT W=0.41u L=40.00n
XX14 net37 nandab VDD VNW PHVT11LL_CKT W=0.41u L=40.00n
XX50 net184 csn net188 VNW PHVT11LL_CKT W=0.295u L=40.00n
XX48 net200 CS net188 VNW PHVT11LL_CKT W=0.205u L=40.00n
XX52 S net188 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX46 orab ci1n net176 VNW PHVT11LL_CKT W=0.42u L=40.00n
XX44 andab CI1 net176 VNW PHVT11LL_CKT W=0.42u L=40.00n
XX54 CO1N net176 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX34 CO0N net152 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX24 orab norab VDD VNW PHVT11LL_CKT W=0.375u L=40.00n
XX30 orab ci0n net152 VNW PHVT11LL_CKT W=0.375u L=40.00n
XX28 andab CI0 net152 VNW PHVT11LL_CKT W=0.375u L=40.00n
XX22 andab nandab VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX18 nandab B VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX15 nandab A VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX2 ci1nnn CI1 VDD VNW PHVT11LL_CKT W=290.00n L=40.00n
XX0 ci0nnn CI0 VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX8 csn CS VDD VNW PHVT11LL_CKT W=290.00n L=40.00n
XX6 ci1n CI1 VDD VNW PHVT11LL_CKT W=290.00n L=40.00n
XX4 ci0n CI0 VDD VNW PHVT11LL_CKT W=290.00n L=40.00n
XX12 norab A net116 VNW PHVT11LL_CKT W=435.00n L=40.00n
XX11 net116 B VDD VNW PHVT11LL_CKT W=435.00n L=40.00n
.ENDS AD2CSCONV2_12TH40
.SUBCKT AD2CSCONV3_12TH40 A B CI0 CI1 CO0N CO1N CS S VDD VSS
XX3 ci1nnn CI1 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX1 ci0nnn CI0 VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX9 csn CS VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX7 ci1n CI1 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX5 ci0n CI0 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX17 net141 B VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX16 nandab A net141 VPW NHVT11LL_CKT W=0.32u L=40.00n
XX31 orab CI0 net152 VPW NHVT11LL_CKT W=0.34u L=40.00n
XX29 andab ci0n net152 VPW NHVT11LL_CKT W=0.34u L=40.00n
XX25 orab norab VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX23 andab nandab VSS VPW NHVT11LL_CKT W=0.325u L=40.00n
XX35 CO0N net152 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX55 CO1N net176 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX47 orab CI1 net176 VPW NHVT11LL_CKT W=0.325u L=40.00n
XX45 andab ci1n net176 VPW NHVT11LL_CKT W=0.325u L=40.00n
XX43 net213 CI1 net184 VPW NHVT11LL_CKT W=0.265u L=40.00n
XX51 net184 CS net188 VPW NHVT11LL_CKT W=0.325u L=40.00n
XX41 net209 ci1nnn net184 VPW NHVT11LL_CKT W=0.34u L=40.00n
XX49 net200 csn net188 VPW NHVT11LL_CKT W=0.325u L=40.00n
XX39 net213 CI0 net200 VPW NHVT11LL_CKT W=0.21u L=40.00n
XX37 net209 ci0nnn net200 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX53 S net188 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX33 net209 net213 VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX27 net213 net37 VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX21 net217 orab VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX20 net37 nandab net217 VPW NHVT11LL_CKT W=0.34u L=40.00n
XX13 norab B VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX10 norab A VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX42 net213 ci1nnn net184 VNW PHVT11LL_CKT W=0.42u L=40.00n
XX40 net209 CI1 net184 VNW PHVT11LL_CKT W=0.42u L=40.00n
XX38 net213 ci0nnn net200 VNW PHVT11LL_CKT W=0.41u L=40.00n
XX36 net209 CI0 net200 VNW PHVT11LL_CKT W=0.41u L=40.00n
XX32 net209 net213 VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX26 net213 net37 VDD VNW PHVT11LL_CKT W=0.41u L=40.00n
XX19 net37 orab VDD VNW PHVT11LL_CKT W=0.41u L=40.00n
XX14 net37 nandab VDD VNW PHVT11LL_CKT W=0.41u L=40.00n
XX50 net184 csn net188 VNW PHVT11LL_CKT W=0.295u L=40.00n
XX48 net200 CS net188 VNW PHVT11LL_CKT W=0.205u L=40.00n
XX52 S net188 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX46 orab ci1n net176 VNW PHVT11LL_CKT W=0.42u L=40.00n
XX44 andab CI1 net176 VNW PHVT11LL_CKT W=0.42u L=40.00n
XX54 CO1N net176 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX34 CO0N net152 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX24 orab norab VDD VNW PHVT11LL_CKT W=0.375u L=40.00n
XX30 orab ci0n net152 VNW PHVT11LL_CKT W=0.375u L=40.00n
XX28 andab CI0 net152 VNW PHVT11LL_CKT W=0.375u L=40.00n
XX22 andab nandab VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX18 nandab B VDD VNW PHVT11LL_CKT W=0.285u L=40.00n
XX15 nandab A VDD VNW PHVT11LL_CKT W=0.285u L=40.00n
XX2 ci1nnn CI1 VDD VNW PHVT11LL_CKT W=290.00n L=40.00n
XX0 ci0nnn CI0 VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX8 csn CS VDD VNW PHVT11LL_CKT W=290.00n L=40.00n
XX6 ci1n CI1 VDD VNW PHVT11LL_CKT W=290.00n L=40.00n
XX4 ci0n CI0 VDD VNW PHVT11LL_CKT W=290.00n L=40.00n
XX12 norab A net116 VNW PHVT11LL_CKT W=0.435u L=40.00n
XX11 net116 B VDD VNW PHVT11LL_CKT W=0.435u L=40.00n
.ENDS AD2CSCONV3_12TH40
.SUBCKT AD2CSCONV4_12TH40 A B CI0 CI1 CO0N CO1N CS S VDD VSS
XX3 ci1nnn CI1 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX1 ci0nnn CI0 VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX9 csn CS VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX7 ci1n CI1 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX5 ci0n CI0 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX17 net141 B VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX16 nandab A net141 VPW NHVT11LL_CKT W=0.32u L=40.00n
XX31 orab CI0 net152 VPW NHVT11LL_CKT W=0.34u L=40.00n
XX29 andab ci0n net152 VPW NHVT11LL_CKT W=0.34u L=40.00n
XX25 orab norab VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX23 andab nandab VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX35 CO0N net152 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX55 CO1N net176 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX47 orab CI1 net176 VPW NHVT11LL_CKT W=0.325u L=40.00n
XX45 andab ci1n net176 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX43 net213 CI1 net184 VPW NHVT11LL_CKT W=0.265u L=40.00n
XX51 net184 CS net188 VPW NHVT11LL_CKT W=0.325u L=40.00n
XX41 net209 ci1nnn net184 VPW NHVT11LL_CKT W=0.315u L=40.00n
XX49 net200 csn net188 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX39 net213 CI0 net200 VPW NHVT11LL_CKT W=0.21u L=40.00n
XX37 net209 ci0nnn net200 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX53 S net188 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX33 net209 net213 VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX27 net213 net37 VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX21 net217 orab VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX20 net37 nandab net217 VPW NHVT11LL_CKT W=0.34u L=40.00n
XX13 norab B VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX10 norab A VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX42 net213 ci1nnn net184 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX40 net209 CI1 net184 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX38 net213 ci0nnn net200 VNW PHVT11LL_CKT W=0.41u L=40.00n
XX36 net209 CI0 net200 VNW PHVT11LL_CKT W=0.41u L=40.00n
XX32 net209 net213 VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX26 net213 net37 VDD VNW PHVT11LL_CKT W=0.41u L=40.00n
XX19 net37 orab VDD VNW PHVT11LL_CKT W=0.41u L=40.00n
XX14 net37 nandab VDD VNW PHVT11LL_CKT W=0.41u L=40.00n
XX50 net184 csn net188 VNW PHVT11LL_CKT W=0.505u L=40.00n
XX48 net200 CS net188 VNW PHVT11LL_CKT W=0.415u L=40.00n
XX52 S net188 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX46 orab ci1n net176 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX44 andab CI1 net176 VNW PHVT11LL_CKT W=0.42u L=40.00n
XX54 CO1N net176 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX34 CO0N net152 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX24 orab norab VDD VNW PHVT11LL_CKT W=0.375u L=40.00n
XX30 orab ci0n net152 VNW PHVT11LL_CKT W=0.375u L=40.00n
XX28 andab CI0 net152 VNW PHVT11LL_CKT W=0.375u L=40.00n
XX22 andab nandab VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX18 nandab B VDD VNW PHVT11LL_CKT W=0.285u L=40.00n
XX15 nandab A VDD VNW PHVT11LL_CKT W=0.285u L=40.00n
XX2 ci1nnn CI1 VDD VNW PHVT11LL_CKT W=0.29u L=40.00n
XX0 ci0nnn CI0 VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX8 csn CS VDD VNW PHVT11LL_CKT W=0.29u L=40.00n
XX6 ci1n CI1 VDD VNW PHVT11LL_CKT W=0.29u L=40.00n
XX4 ci0n CI0 VDD VNW PHVT11LL_CKT W=0.29u L=40.00n
XX12 norab A net116 VNW PHVT11LL_CKT W=0.435u L=40.00n
XX11 net116 B VDD VNW PHVT11LL_CKT W=0.435u L=40.00n
.ENDS AD2CSCONV4_12TH40
.SUBCKT ADH1CINV2C_12TH40 A CIN CO S VDD VSS
XX7 net_65 acinn net_33 VPW NHVT11LL_CKT W=465.00n L=40.00n
XX13 S net_65 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX11 net_13 net35 VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX1 net35 CIN VSS VPW NHVT11LL_CKT W=300.00n L=40.00n
XX10 acinn A net_13 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX15 CO acinn VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX8 net_33 net35 VSS VPW NHVT11LL_CKT W=465.00n L=40.00n
XX4 net_33 A VSS VPW NHVT11LL_CKT W=465.00n L=40.00n
XX6 net_65 acinn VDD VNW PHVT11LL_CKT W=305.00n L=40.00n
XX5 acinn A VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX9 acinn net35 VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX12 S net_65 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX2 net_68 net35 VDD VNW PHVT11LL_CKT W=565.00n L=40.00n
XX14 CO acinn VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX0 net35 CIN VDD VNW PHVT11LL_CKT W=340.00n L=40.00n
XX3 net_65 A net_68 VNW PHVT11LL_CKT W=565.00n L=40.00n
.ENDS ADH1CINV2C_12TH40
.SUBCKT ADH1CINV2_12TH40 A CIN CO S VDD VSS
XX15 net45 CIN S VPW NHVT11LL_CKT W=540.00n L=40.00n
XX14 net46 net35 S VPW NHVT11LL_CKT W=540.00n L=40.00n
XX13 CO net_53 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX12 net_17 net35 VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX11 net_53 A net_17 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX10 net35 CIN VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX9 net45 net46 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX8 net46 A VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX7 net45 net35 S VNW PHVT11LL_CKT W=610.00n L=40.00n
XX6 net46 CIN S VNW PHVT11LL_CKT W=610.00n L=40.00n
XX5 CO net_53 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX4 net_53 net35 VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX3 net_53 A VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX2 net35 CIN VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
XX1 net45 net46 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX0 net46 A VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
.ENDS ADH1CINV2_12TH40
.SUBCKT ADH1CINV3C_12TH40 A CIN CO S VDD VSS
XX7 net_65 acinn net_33 VPW NHVT11LL_CKT W=540.00n L=40.00n
XX13 S net_65 VSS VPW NHVT11LL_CKT W=0.78u L=40.00n
XX11 net_13 net35 VSS VPW NHVT11LL_CKT W=450.00n L=40.00n
XX1 net35 CIN VSS VPW NHVT11LL_CKT W=420.00n L=40.00n
XX10 acinn A net_13 VPW NHVT11LL_CKT W=450.00n L=40.00n
XX15 CO acinn VSS VPW NHVT11LL_CKT W=0.78u L=40.00n
XX8 net_33 net35 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX4 net_33 A VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX6 net_65 acinn VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX5 acinn A VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX9 acinn net35 VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX12 S net_65 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX2 net_68 net35 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX14 CO acinn VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX0 net35 CIN VDD VNW PHVT11LL_CKT W=480.00n L=40.00n
XX3 net_65 A net_68 VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS ADH1CINV3C_12TH40
.SUBCKT ADH1CINV3_12TH40 A CIN CO S VDD VSS
XX15 net45 CIN S VPW NHVT11LL_CKT W=760.00n L=40.00n
XX14 net46 net35 S VPW NHVT11LL_CKT W=760.00n L=40.00n
XX13 CO net_53 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX12 net_17 net35 VSS VPW NHVT11LL_CKT W=450.00n L=40.00n
XX11 net_53 A net_17 VPW NHVT11LL_CKT W=450.00n L=40.00n
XX10 net35 CIN VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX9 net45 net46 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX8 net46 A VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX7 net45 net35 S VNW PHVT11LL_CKT W=860.00n L=40.00n
XX6 net46 CIN S VNW PHVT11LL_CKT W=860.00n L=40.00n
XX5 CO net_53 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX4 net_53 net35 VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX3 net_53 A VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX2 net35 CIN VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX1 net45 net46 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX0 net46 A VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS ADH1CINV3_12TH40
.SUBCKT ADH1CINV4C_12TH40 A CIN CO S VDD VSS
XX6 net_64 acinn VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX5 acinn A VDD VNW PHVT11LL_CKT W=550.00n L=40.00n
XX9 acinn net35 VDD VNW PHVT11LL_CKT W=550.00n L=40.00n
XX12 S net_64 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX2 net_67 net35 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX14 CO acinn VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 net35 CIN VDD VNW PHVT11LL_CKT W=480.00n L=40.00n
XX3 net_64 A net_67 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX7 net_64 acinn net_96 VPW NHVT11LL_CKT W=540.00n L=40.00n
XX13 S net_64 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX11 net_116 net35 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX1 net35 CIN VSS VPW NHVT11LL_CKT W=420.00n L=40.00n
XX10 acinn A net_116 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX15 CO acinn VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX8 net_96 net35 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX4 net_96 A VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
.ENDS ADH1CINV4C_12TH40
.SUBCKT ADH1CINV4_12TH40 A CIN CO S VDD VSS
XX15 net45 CIN S VPW NHVT11LL_CKT W=1.08u L=40.00n
XX14 net46 net35 S VPW NHVT11LL_CKT W=1.08u L=40.00n
XX13 CO net_53 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX12 net_17 net35 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX11 net_53 A net_17 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX10 net35 CIN VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX9 net45 net46 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX8 net46 A VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX7 net45 net35 S VNW PHVT11LL_CKT W=1.22u L=40.00n
XX6 net46 CIN S VNW PHVT11LL_CKT W=1.22u L=40.00n
XX5 CO net_53 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX4 net_53 net35 VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX3 net_53 A VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX2 net35 CIN VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 net45 net46 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 net46 A VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS ADH1CINV4_12TH40
.SUBCKT ADH1CONV2_12TH40 A CI CON S VDD VSS
XX6 net45 net35 S VPW NHVT11LL_CKT W=540.00n L=40.00n
XX5 net46 CI S VPW NHVT11LL_CKT W=540.00n L=40.00n
XX4 net_41 CI VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX3 CON A net_41 VPW NHVT11LL_CKT W=540.00n L=40.00n
XX2 net35 CI VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX1 net45 net46 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX0 net46 A VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX13 net45 CI S VNW PHVT11LL_CKT W=610.00n L=40.00n
XX12 net46 net35 S VNW PHVT11LL_CKT W=610.00n L=40.00n
XX11 CON CI VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX10 CON A VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX9 net35 CI VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
XX8 net45 net46 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX7 net46 A VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
.ENDS ADH1CONV2_12TH40
.SUBCKT ADH1CONV3_12TH40 A CI CON S VDD VSS
XX6 net45 net35 S VPW NHVT11LL_CKT W=760.00n L=40.00n
XX5 net46 CI S VPW NHVT11LL_CKT W=760.00n L=40.00n
XX4 net_41 CI VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX3 CON A net_41 VPW NHVT11LL_CKT W=760.00n L=40.00n
XX2 net35 CI VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX1 net45 net46 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX0 net46 A VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX13 net45 CI S VNW PHVT11LL_CKT W=860.00n L=40.00n
XX12 net46 net35 S VNW PHVT11LL_CKT W=860.00n L=40.00n
XX11 CON CI VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX10 CON A VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX9 net35 CI VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX8 net45 net46 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX7 net46 A VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS ADH1CONV3_12TH40
.SUBCKT ADH1CONV4_12TH40 A CI CON S VDD VSS
XX6 net45 net35 S VPW NHVT11LL_CKT W=1.08u L=40.00n
XX5 net46 CI S VPW NHVT11LL_CKT W=1.08u L=40.00n
XX4 net_41 CI VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX3 CON A net_41 VPW NHVT11LL_CKT W=1.08u L=40.00n
XX2 net35 CI VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX1 net45 net46 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX0 net46 A VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX13 net45 CI S VNW PHVT11LL_CKT W=1.22u L=40.00n
XX12 net46 net35 S VNW PHVT11LL_CKT W=1.22u L=40.00n
XX11 CON CI VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX10 CON A VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX9 net35 CI VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX8 net45 net46 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX7 net46 A VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS ADH1CONV4_12TH40
.SUBCKT ADH1CSCINV2_12TH40 A CIN CO CS S VDD VSS
XX20 S net17 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX13 an csn net17 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX15 net34 CS net17 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX11 an CIN net34 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX21 CO CIN VSS VPW NHVT11LL_CKT W=275.00n L=40.00n
XX18 CO an VSS VPW NHVT11LL_CKT W=275.00n L=40.00n
XX9 net30 an VSS VPW NHVT11LL_CKT W=340.00n L=40.00n
XX8 net34 cinn net30 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX5 csn CS VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX3 cinn CIN VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX1 an A VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX10 an cinn net34 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX14 net34 csn net17 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX12 an CS net17 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX19 S net17 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX17 CO CIN net69 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX16 net69 an VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX7 net34 CIN net77 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX6 net77 an VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX4 csn CS VDD VNW PHVT11LL_CKT W=290.00n L=40.00n
XX2 cinn CIN VDD VNW PHVT11LL_CKT W=290.00n L=40.00n
XX0 an A VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS ADH1CSCINV2_12TH40
.SUBCKT ADH1CSCINV3_12TH40 A CIN CO CS S VDD VSS
XX20 S net17 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX13 an csn net17 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX15 net34 CS net17 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX11 an CIN net34 VPW NHVT11LL_CKT W=395.00n L=40.00n
XX21 CO CIN VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX18 CO an VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX9 net30 an VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX8 net34 cinn net30 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX5 csn CS VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX3 cinn CIN VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX1 an A VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX10 an cinn net34 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX14 net34 csn net17 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX12 an CS net17 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX19 S net17 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX17 CO CIN net69 VNW PHVT11LL_CKT W=860.00n L=40.00n
XX16 net69 an VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX7 net34 CIN net77 VNW PHVT11LL_CKT W=460.00n L=40.00n
XX6 net77 an VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
XX4 csn CS VDD VNW PHVT11LL_CKT W=330.00n L=40.00n
XX2 cinn CIN VDD VNW PHVT11LL_CKT W=330.00n L=40.00n
XX0 an A VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS ADH1CSCINV3_12TH40
.SUBCKT ADH1CSCINV4_12TH40 A CIN CO CS S VDD VSS
XX20 S net17 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX13 an csn net17 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX15 net34 CS net17 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX11 an CIN net34 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX21 CO CIN VSS VPW NHVT11LL_CKT W=550.00n L=40.00n
XX18 CO an VSS VPW NHVT11LL_CKT W=550.00n L=40.00n
XX9 net30 an VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX8 net34 cinn net30 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX5 csn CS VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX3 cinn CIN VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX1 an A VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX10 an cinn net34 VNW PHVT11LL_CKT W=500.0n L=40.00n
XX14 net34 csn net17 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX12 an CS net17 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX19 S net17 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX17 CO CIN net69 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX16 net69 an VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX7 net34 CIN net77 VNW PHVT11LL_CKT W=460.00n L=40.00n
XX6 net77 an VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
XX4 csn CS VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
XX2 cinn CIN VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
XX0 an A VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS ADH1CSCINV4_12TH40
.SUBCKT ADH1CSCONV2_12TH40 A CI CON CS S VDD VSS
XX11 an cin net78 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX15 net78 CS net57 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX13 an csn net57 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX21 S net57 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX19 net66 A VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX18 CON CI net66 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX9 net74 an VSS VPW NHVT11LL_CKT W=340.00n L=40.00n
XX8 net78 CI net74 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX5 csn CS VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX3 cin CI VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX1 an A VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX10 an CI net78 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX14 net78 csn net57 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX12 an CS net57 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX20 S net57 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX17 CON CI VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX16 CON A VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX7 net78 cin net33 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX6 net33 an VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX4 csn CS VDD VNW PHVT11LL_CKT W=290.00n L=40.00n
XX2 cin CI VDD VNW PHVT11LL_CKT W=290.00n L=40.00n
XX0 an A VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS ADH1CSCONV2_12TH40
.SUBCKT ADH1CSCONV3_12TH40 A CI CON CS S VDD VSS
XX11 an cin net78 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX15 net78 CS net57 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX13 an csn net57 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX21 S net57 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX19 net66 A VSS VPW NHVT11LL_CKT W=860.00n L=40.00n
XX18 CON CI net66 VPW NHVT11LL_CKT W=860.00n L=40.00n
XX9 net74 an VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX8 net78 CI net74 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX5 csn CS VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX3 cin CI VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX1 an A VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX10 an CI net78 VNW PHVT11LL_CKT W=0.45u L=40.00n
XX14 net78 csn net57 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX12 an CS net57 VNW PHVT11LL_CKT W=0.54u L=40.00n
XX20 S net57 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX17 CON CI VDD VNW PHVT11LL_CKT W=760.00n L=40.00n
XX16 CON A VDD VNW PHVT11LL_CKT W=760.00n L=40.00n
XX7 net78 cin net33 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX6 net33 an VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
XX4 csn CS VDD VNW PHVT11LL_CKT W=330.00n L=40.00n
XX2 cin CI VDD VNW PHVT11LL_CKT W=330.00n L=40.00n
XX0 an A VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
.ENDS ADH1CSCONV3_12TH40
.SUBCKT ADH1CSCONV4_12TH40 A CI CON CS S VDD VSS
XX11 an cin net78 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX15 net78 CS net57 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX13 an csn net57 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX21 S net57 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX19 net66 A VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX18 CON CI net66 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX9 net74 an VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX8 net78 CI net74 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX5 csn CS VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX3 cin CI VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX1 an A VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX10 an CI net78 VNW PHVT11LL_CKT W=0.45u L=40.00n
XX14 net78 csn net57 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX12 an CS net57 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX20 S net57 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX17 CON CI VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX16 CON A VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX7 net78 cin net33 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX6 net33 an VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX4 csn CS VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
XX2 cin CI VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
XX0 an A VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS ADH1CSCONV4_12TH40
.SUBCKT ADH1V2C_12TH40 A B CO S VDD VSS
XX11 S net17 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX10 net17 nandab net9 VPW NHVT11LL_CKT W=300.00n L=40.00n
XX29 net9 A VSS VPW NHVT11LL_CKT W=300.00n L=40.00n
XX2 net9 B VSS VPW NHVT11LL_CKT W=300.00n L=40.00n
XX4 CO nandab VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX8 net25 B VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX9 nandab A net25 VPW NHVT11LL_CKT W=500.00n L=40.00n
XX3 S net17 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 net17 nandab VDD VNW PHVT11LL_CKT W=195.00n L=40.00n
XX6 net48 B VDD VNW PHVT11LL_CKT W=360.00n L=40.00n
XX7 net17 A net48 VNW PHVT11LL_CKT W=360.00n L=40.00n
XX5 CO nandab VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX28 nandab A VDD VNW PHVT11LL_CKT W=330.00n L=40.00n
XX0 nandab B VDD VNW PHVT11LL_CKT W=330.00n L=40.00n
.ENDS ADH1V2C_12TH40
.SUBCKT ADH1V2_12TH40 A B CO S VDD VSS
XX14 net5 A VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX13 net41 B net5 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX17 CO net41 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX7 net37 bn net20 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX9 net33 B net20 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX1 bn B VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX11 S net20 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX5 net33 net37 VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX3 net37 A VSS VPW NHVT11LL_CKT W=430.00n L=40.00n
XX12 net41 A VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX8 net33 bn net20 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX15 net41 B VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX4 net33 net37 VDD VNW PHVT11LL_CKT W=390.00n L=40.00n
XX10 S net20 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX16 CO net41 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX0 bn B VDD VNW PHVT11LL_CKT W=290.00n L=40.00n
XX6 net37 B net20 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX2 net37 A VDD VNW PHVT11LL_CKT W=520.00n L=40.00n
.ENDS ADH1V2_12TH40
.SUBCKT ADH1V3C_12TH40 A B CO S VDD VSS
XX11 S net17 VSS VPW NHVT11LL_CKT W=0.75u L=40.00n
XX10 net17 nandab net9 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX29 net9 A VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX2 net9 B VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX4 CO nandab VSS VPW NHVT11LL_CKT W=0.75u L=40.00n
XX8 net25 B VSS VPW NHVT11LL_CKT W=0.575u L=40.00n
XX9 nandab A net25 VPW NHVT11LL_CKT W=0.575u L=40.00n
XX3 S net17 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX1 net17 nandab VDD VNW PHVT11LL_CKT W=0.26u L=40.00n
XX6 net48 B VDD VNW PHVT11LL_CKT W=0.485u L=40.00n
XX7 net17 A net48 VNW PHVT11LL_CKT W=0.485u L=40.00n
XX5 CO nandab VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX28 nandab A VDD VNW PHVT11LL_CKT W=0.375u L=40.00n
XX0 nandab B VDD VNW PHVT11LL_CKT W=0.375u L=40.00n
.ENDS ADH1V3C_12TH40
.SUBCKT ADH1V3_12TH40 A B CO S VDD VSS
XX14 net5 A VSS VPW NHVT11LL_CKT W=450.00n L=40.00n
XX13 net41 B net5 VPW NHVT11LL_CKT W=450.00n L=40.00n
XX17 CO net41 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX7 net37 bn net20 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX9 net33 B net20 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX1 bn B VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX11 S net20 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX5 net33 net37 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX3 net37 A VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX12 net41 A VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX8 net33 bn net20 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX15 net41 B VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX4 net33 net37 VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX10 S net20 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX16 CO net41 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX0 bn B VDD VNW PHVT11LL_CKT W=330.00n L=40.00n
XX6 net37 B net20 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX2 net37 A VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
.ENDS ADH1V3_12TH40
.SUBCKT ADH1V4C_12TH40 A B CO S VDD VSS
XX11 S net17 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX10 net17 nandab net9 VPW NHVT11LL_CKT W=0.505u L=40.00n
XX29 net9 A VSS VPW NHVT11LL_CKT W=0.505u L=40.00n
XX2 net9 B VSS VPW NHVT11LL_CKT W=0.505u L=40.00n
XX4 CO nandab VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX8 net25 B VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX9 nandab A net25 VPW NHVT11LL_CKT W=0.61u L=40.00n
XX3 S net17 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 net17 nandab VDD VNW PHVT11LL_CKT W=0.325u L=40.00n
XX6 net48 B VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX7 net17 A net48 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX5 CO nandab VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX28 nandab A VDD VNW PHVT11LL_CKT W=0.395u L=40.00n
XX0 nandab B VDD VNW PHVT11LL_CKT W=0.395u L=40.00n
.ENDS ADH1V4C_12TH40
.SUBCKT ADH1V4_12TH40 A B CO S VDD VSS
XX14 net5 A VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX13 net41 B net5 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX17 CO net41 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX7 net37 bn net20 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX9 net33 B net20 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX1 bn B VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX11 S net20 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX5 net33 net37 VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX3 net37 A VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX12 net41 A VDD VNW PHVT11LL_CKT W=550.00n L=40.00n
XX8 net33 bn net20 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX15 net41 B VDD VNW PHVT11LL_CKT W=550.00n L=40.00n
XX4 net33 net37 VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
XX10 S net20 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX16 CO net41 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 bn B VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX6 net37 B net20 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX2 net37 A VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS ADH1V4_12TH40
.SUBCKT AND2V0_12TH40 A1 A2 Z VDD VSS
XX6 Z net037 VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX9 net037 A1 net16 VPW NHVT11LL_CKT W=165.00n L=40.00n
XX8 net16 A2 VSS VPW NHVT11LL_CKT W=165.00n L=40.00n
XX0 net037 A2 VDD VNW PHVT11LL_CKT W=145.00n L=40.00n
XX28 net037 A1 VDD VNW PHVT11LL_CKT W=145.00n L=40.00n
XX5 Z net037 VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
.ENDS AND2V0_12TH40
.SUBCKT AND2V10RD_12TH40 A1 A2 Z VDD VSS
XX6 Z net037 VSS VPW NHVT11LL_CKT W=2.7u L=40.00n
XX9 net037 A1 net16 VPW NHVT11LL_CKT W=3.05u L=40.00n
XX8 net16 A2 VSS VPW NHVT11LL_CKT W=3.05u L=40.00n
XX0 net037 A2 VDD VNW PHVT11LL_CKT W=2.00u L=40.00n
XX28 net037 A1 VDD VNW PHVT11LL_CKT W=2.00u L=40.00n
XX5 Z net037 VDD VNW PHVT11LL_CKT W=3.05u L=40.00n
.ENDS AND2V10RD_12TH40
.SUBCKT AND2V12_12TH40 A1 A2 Z VDD VSS
XX6 Z net037 VSS VPW NHVT11LL_CKT W=3.24u L=40.00n
XX9 net037 A1 net16 VPW NHVT11LL_CKT W=1.71u L=40.00n
XX8 net16 A2 VSS VPW NHVT11LL_CKT W=1.71u L=40.00n
XX0 net037 A2 VDD VNW PHVT11LL_CKT W=1.53u L=40.00n
XX28 net037 A1 VDD VNW PHVT11LL_CKT W=1.53u L=40.00n
XX5 Z net037 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
.ENDS AND2V12_12TH40
.SUBCKT AND2V16_12TH40 A1 A2 Z VDD VSS
XX6 Z net037 VSS VPW NHVT11LL_CKT W=4.32u L=40.00n
XX9 net037 A1 net16 VPW NHVT11LL_CKT W=2.3u L=40.00n
XX8 net16 A2 VSS VPW NHVT11LL_CKT W=2.3u L=40.00n
XX0 net037 A2 VDD VNW PHVT11LL_CKT W=2.08u L=40.00n
XX28 net037 A1 VDD VNW PHVT11LL_CKT W=2.08u L=40.00n
XX5 Z net037 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
.ENDS AND2V16_12TH40
.SUBCKT AND2V1RD_12TH40 A1 A2 Z VDD VSS
XX6 Z net037 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX9 net037 A1 net16 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX8 net16 A2 VSS VPW NHVT11LL_CKT W=430.00n L=40.00n
XX0 net037 A2 VDD VNW PHVT11LL_CKT W=280.00n L=40.00n
XX28 net037 A1 VDD VNW PHVT11LL_CKT W=280.00n L=40.00n
XX5 Z net037 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
.ENDS AND2V1RD_12TH40
.SUBCKT AND2V1_12TH40 A1 A2 Z VDD VSS
XX6 Z net037 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX9 net037 A1 net16 VPW NHVT11LL_CKT W=225.00n L=40.00n
XX8 net16 A2 VSS VPW NHVT11LL_CKT W=225.00n L=40.00n
XX0 net037 A2 VDD VNW PHVT11LL_CKT W=200.00n L=40.00n
XX28 net037 A1 VDD VNW PHVT11LL_CKT W=200.00n L=40.00n
XX5 Z net037 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
.ENDS AND2V1_12TH40
.SUBCKT AND2V20_12TH40 A1 A2 Z VDD VSS
XX6 Z net037 VSS VPW NHVT11LL_CKT W=5.4u L=40.00n
XX9 net037 A1 net16 VPW NHVT11LL_CKT W=3.05u L=40.00n
XX8 net16 A2 VSS VPW NHVT11LL_CKT W=3.05u L=40.00n
XX0 net037 A2 VDD VNW PHVT11LL_CKT W=2.75u L=40.00n
XX28 net037 A1 VDD VNW PHVT11LL_CKT W=2.75u L=40.00n
XX5 Z net037 VDD VNW PHVT11LL_CKT W=6.1u L=40.00n
.ENDS AND2V20_12TH40
.SUBCKT AND2V24_12TH40 A1 A2 Z VDD VSS
XX6 Z net037 VSS VPW NHVT11LL_CKT W=6.48u L=40.00n
XX9 net037 A1 net16 VPW NHVT11LL_CKT W=3.66u L=40.00n
XX8 net16 A2 VSS VPW NHVT11LL_CKT W=3.66u L=40.00n
XX0 net037 A2 VDD VNW PHVT11LL_CKT W=3.3u L=40.00n
XX28 net037 A1 VDD VNW PHVT11LL_CKT W=3.3u L=40.00n
XX5 Z net037 VDD VNW PHVT11LL_CKT W=7.32u L=40.00n
.ENDS AND2V24_12TH40
.SUBCKT AND2V2RD_12TH40 A1 A2 Z VDD VSS
XX6 Z net037 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX9 net037 A1 net16 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX8 net16 A2 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX0 net037 A2 VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX28 net037 A1 VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX5 Z net037 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS AND2V2RD_12TH40
.SUBCKT AND2V2_12TH40 A1 A2 Z VDD VSS
XX6 Z net037 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX9 net037 A1 net16 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX8 net16 A2 VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX0 net037 A2 VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX28 net037 A1 VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX5 Z net037 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS AND2V2_12TH40
.SUBCKT AND2V3_12TH40 A1 A2 Z VDD VSS
XX6 Z net037 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX9 net037 A1 net16 VPW NHVT11LL_CKT W=450.00n L=40.00n
XX8 net16 A2 VSS VPW NHVT11LL_CKT W=450.00n L=40.00n
XX0 net037 A2 VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX28 net037 A1 VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX5 Z net037 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
.ENDS AND2V3_12TH40
.SUBCKT AND2V4RD_12TH40 A1 A2 Z VDD VSS
XX6 Z net037 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX9 net037 A1 net16 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX8 net16 A2 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX0 net037 A2 VDD VNW PHVT11LL_CKT W=800.00n L=40.00n
XX28 net037 A1 VDD VNW PHVT11LL_CKT W=800.00n L=40.00n
XX5 Z net037 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS AND2V4RD_12TH40
.SUBCKT AND2V4_12TH40 A1 A2 Z VDD VSS
XX6 Z net037 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX9 net037 A1 net16 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX8 net16 A2 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX0 net037 A2 VDD VNW PHVT11LL_CKT W=550.00n L=40.00n
XX28 net037 A1 VDD VNW PHVT11LL_CKT W=550.00n L=40.00n
XX5 Z net037 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS AND2V4_12TH40
.SUBCKT AND2V6RD_12TH40 A1 A2 Z VDD VSS
XX6 Z net037 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX9 net037 A1 net16 VPW NHVT11LL_CKT W=1.845u L=40.00n
XX8 net16 A2 VSS VPW NHVT11LL_CKT W=1.845u L=40.00n
XX0 net037 A2 VDD VNW PHVT11LL_CKT W=1.2u L=40.00n
XX28 net037 A1 VDD VNW PHVT11LL_CKT W=1.2u L=40.00n
XX5 Z net037 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS AND2V6RD_12TH40
.SUBCKT AND2V6_12TH40 A1 A2 Z VDD VSS
XX6 Z net037 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX9 net037 A1 net16 VPW NHVT11LL_CKT W=860.00n L=40.00n
XX8 net16 A2 VSS VPW NHVT11LL_CKT W=860.00n L=40.00n
XX0 net037 A2 VDD VNW PHVT11LL_CKT W=780.00n L=40.00n
XX28 net037 A1 VDD VNW PHVT11LL_CKT W=780.00n L=40.00n
XX5 Z net037 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS AND2V6_12TH40
.SUBCKT AND2V8RD_12TH40 A1 A2 Z VDD VSS
XX6 Z net037 VSS VPW NHVT11LL_CKT W=2.14u L=40.00n
XX9 net037 A1 net16 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX8 net16 A2 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX0 net037 A2 VDD VNW PHVT11LL_CKT W=1.6u L=40.00n
XX28 net037 A1 VDD VNW PHVT11LL_CKT W=1.6u L=40.00n
XX5 Z net037 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS AND2V8RD_12TH40
.SUBCKT AND2V8_12TH40 A1 A2 Z VDD VSS
XX6 Z net037 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX9 net037 A1 net16 VPW NHVT11LL_CKT W=1.08u L=40.00n
XX8 net16 A2 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX0 net037 A2 VDD VNW PHVT11LL_CKT W=960.00n L=40.00n
XX28 net037 A1 VDD VNW PHVT11LL_CKT W=960.00n L=40.00n
XX5 Z net037 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS AND2V8_12TH40
.SUBCKT AND3V0_12TH40 A1 A2 A3 Z VDD VSS
XX6 Z net053 VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX2 net053 A1 net17 VPW NHVT11LL_CKT W=380.00n L=40.00n
XX9 net17 A2 net21 VPW NHVT11LL_CKT W=380.00n L=40.00n
XX8 net21 A3 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX1 net053 A3 VDD VNW PHVT11LL_CKT W=225.00n L=40.00n
XX0 net053 A2 VDD VNW PHVT11LL_CKT W=225.00n L=40.00n
XX28 net053 A1 VDD VNW PHVT11LL_CKT W=225.00n L=40.00n
XX5 Z net053 VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
.ENDS AND3V0_12TH40
.SUBCKT AND3V10RD_12TH40 A1 A2 A3 Z VDD VSS
XX6 Z net053 VSS VPW NHVT11LL_CKT W=2.7u L=40.00n
XX2 net053 A1 net17 VPW NHVT11LL_CKT W=3.99u L=40.00n
XX9 net17 A2 net21 VPW NHVT11LL_CKT W=3.99u L=40.00n
XX8 net21 A3 VSS VPW NHVT11LL_CKT W=3.99u L=40.00n
XX1 net053 A3 VDD VNW PHVT11LL_CKT W=2.03u L=40.00n
XX0 net053 A2 VDD VNW PHVT11LL_CKT W=2.03u L=40.00n
XX28 net053 A1 VDD VNW PHVT11LL_CKT W=2.03u L=40.00n
XX5 Z net053 VDD VNW PHVT11LL_CKT W=3.05u L=40.00n
.ENDS AND3V10RD_12TH40
.SUBCKT AND3V12_12TH40 A1 A2 A3 Z VDD VSS
XX6 Z net053 VSS VPW NHVT11LL_CKT W=3.24u L=40.00n
XX2 net053 A1 net17 VPW NHVT11LL_CKT W=3.24u L=40.00n
XX9 net17 A2 net21 VPW NHVT11LL_CKT W=3.24u L=40.00n
XX8 net21 A3 VSS VPW NHVT11LL_CKT W=3.24u L=40.00n
XX1 net053 A3 VDD VNW PHVT11LL_CKT W=1.95u L=40.00n
XX0 net053 A2 VDD VNW PHVT11LL_CKT W=1.95u L=40.00n
XX28 net053 A1 VDD VNW PHVT11LL_CKT W=1.95u L=40.00n
XX5 Z net053 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
.ENDS AND3V12_12TH40
.SUBCKT AND3V16_12TH40 A1 A2 A3 Z VDD VSS
XX6 Z net053 VSS VPW NHVT11LL_CKT W=4.32u L=40.00n
XX2 net053 A1 net17 VPW NHVT11LL_CKT W=4.32u L=40.00n
XX9 net17 A2 net21 VPW NHVT11LL_CKT W=4.32u L=40.00n
XX8 net21 A3 VSS VPW NHVT11LL_CKT W=4.32u L=40.00n
XX1 net053 A3 VDD VNW PHVT11LL_CKT W=2.6u L=40.00n
XX0 net053 A2 VDD VNW PHVT11LL_CKT W=2.6u L=40.00n
XX28 net053 A1 VDD VNW PHVT11LL_CKT W=2.6u L=40.00n
XX5 Z net053 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
.ENDS AND3V16_12TH40
.SUBCKT AND3V1RD_12TH40 A1 A2 A3 Z VDD VSS
XX6 Z net053 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX2 net053 A1 net17 VPW NHVT11LL_CKT W=560.00n L=40.00n
XX9 net17 A2 net21 VPW NHVT11LL_CKT W=560.00n L=40.00n
XX8 net21 A3 VSS VPW NHVT11LL_CKT W=560.00n L=40.00n
XX1 net053 A3 VDD VNW PHVT11LL_CKT W=280.00n L=40.00n
XX0 net053 A2 VDD VNW PHVT11LL_CKT W=280.00n L=40.00n
XX28 net053 A1 VDD VNW PHVT11LL_CKT W=280.00n L=40.00n
XX5 Z net053 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
.ENDS AND3V1RD_12TH40
.SUBCKT AND3V1_12TH40 A1 A2 A3 Z VDD VSS
XX6 Z net053 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX2 net053 A1 net17 VPW NHVT11LL_CKT W=460.00n L=40.00n
XX9 net17 A2 net21 VPW NHVT11LL_CKT W=460.00n L=40.00n
XX8 net21 A3 VSS VPW NHVT11LL_CKT W=460.00n L=40.00n
XX1 net053 A3 VDD VNW PHVT11LL_CKT W=275.00n L=40.00n
XX0 net053 A2 VDD VNW PHVT11LL_CKT W=275.00n L=40.00n
XX28 net053 A1 VDD VNW PHVT11LL_CKT W=275.00n L=40.00n
XX5 Z net053 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
.ENDS AND3V1_12TH40
.SUBCKT AND3V2RD_12TH40 A1 A2 A3 Z VDD VSS
XX6 Z net053 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX2 net053 A1 net17 VPW NHVT11LL_CKT W=800.00n L=40.00n
XX9 net17 A2 net21 VPW NHVT11LL_CKT W=800.00n L=40.00n
XX8 net21 A3 VSS VPW NHVT11LL_CKT W=800.00n L=40.00n
XX1 net053 A3 VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX0 net053 A2 VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX28 net053 A1 VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX5 Z net053 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS AND3V2RD_12TH40
.SUBCKT AND3V2_12TH40 A1 A2 A3 Z VDD VSS
XX6 Z net053 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX2 net053 A1 net17 VPW NHVT11LL_CKT W=540.00n L=40.00n
XX9 net17 A2 net21 VPW NHVT11LL_CKT W=540.00n L=40.00n
XX8 net21 A3 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX1 net053 A3 VDD VNW PHVT11LL_CKT W=325.00n L=40.00n
XX0 net053 A2 VDD VNW PHVT11LL_CKT W=325.00n L=40.00n
XX28 net053 A1 VDD VNW PHVT11LL_CKT W=325.00n L=40.00n
XX5 Z net053 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS AND3V2_12TH40
.SUBCKT AND3V3_12TH40 A1 A2 A3 Z VDD VSS
XX6 Z net053 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX2 net053 A1 net17 VPW NHVT11LL_CKT W=590.00n L=40.00n
XX9 net17 A2 net21 VPW NHVT11LL_CKT W=590.00n L=40.00n
XX8 net21 A3 VSS VPW NHVT11LL_CKT W=590.00n L=40.00n
XX1 net053 A3 VDD VNW PHVT11LL_CKT W=275.00n L=40.00n
XX0 net053 A2 VDD VNW PHVT11LL_CKT W=275.00n L=40.00n
XX28 net053 A1 VDD VNW PHVT11LL_CKT W=275.00n L=40.00n
XX5 Z net053 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS AND3V3_12TH40
.SUBCKT AND3V4RD_12TH40 A1 A2 A3 Z VDD VSS
XX6 Z net053 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX2 net053 A1 net17 VPW NHVT11LL_CKT W=1.59u L=40.00n
XX9 net17 A2 net21 VPW NHVT11LL_CKT W=1.59u L=40.00n
XX8 net21 A3 VSS VPW NHVT11LL_CKT W=1.59u L=40.00n
XX1 net053 A3 VDD VNW PHVT11LL_CKT W=810.00n L=40.00n
XX0 net053 A2 VDD VNW PHVT11LL_CKT W=810.00n L=40.00n
XX28 net053 A1 VDD VNW PHVT11LL_CKT W=810.00n L=40.00n
XX5 Z net053 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS AND3V4RD_12TH40
.SUBCKT AND3V4_12TH40 A1 A2 A3 Z VDD VSS
XX6 Z net053 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX2 net053 A1 net17 VPW NHVT11LL_CKT W=1.08u L=40.00n
XX9 net17 A2 net21 VPW NHVT11LL_CKT W=1.08u L=40.00n
XX8 net21 A3 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX1 net053 A3 VDD VNW PHVT11LL_CKT W=650.00n L=40.00n
XX0 net053 A2 VDD VNW PHVT11LL_CKT W=650.00n L=40.00n
XX28 net053 A1 VDD VNW PHVT11LL_CKT W=650.00n L=40.00n
XX5 Z net053 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS AND3V4_12TH40
.SUBCKT AND3V6RD_12TH40 A1 A2 A3 Z VDD VSS
XX6 Z net053 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX2 net053 A1 net17 VPW NHVT11LL_CKT W=2.4u L=40.00n
XX9 net17 A2 net21 VPW NHVT11LL_CKT W=2.4u L=40.00n
XX8 net21 A3 VSS VPW NHVT11LL_CKT W=2.4u L=40.00n
XX1 net053 A3 VDD VNW PHVT11LL_CKT W=1.2u L=40.00n
XX0 net053 A2 VDD VNW PHVT11LL_CKT W=1.2u L=40.00n
XX28 net053 A1 VDD VNW PHVT11LL_CKT W=1.2u L=40.00n
XX5 Z net053 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS AND3V6RD_12TH40
.SUBCKT AND3V6_12TH40 A1 A2 A3 Z VDD VSS
XX6 Z net053 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX2 net053 A1 net17 VPW NHVT11LL_CKT W=1.62u L=40.00n
XX9 net17 A2 net21 VPW NHVT11LL_CKT W=1.62u L=40.00n
XX8 net21 A3 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX1 net053 A3 VDD VNW PHVT11LL_CKT W=975.00n L=40.00n
XX0 net053 A2 VDD VNW PHVT11LL_CKT W=975.00n L=40.00n
XX28 net053 A1 VDD VNW PHVT11LL_CKT W=975.00n L=40.00n
XX5 Z net053 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS AND3V6_12TH40
.SUBCKT AND3V8RD_12TH40 A1 A2 A3 Z VDD VSS
XX6 Z net053 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX2 net053 A1 net17 VPW NHVT11LL_CKT W=3.18u L=40.00n
XX9 net17 A2 net21 VPW NHVT11LL_CKT W=3.18u L=40.00n
XX8 net21 A3 VSS VPW NHVT11LL_CKT W=3.18u L=40.00n
XX1 net053 A3 VDD VNW PHVT11LL_CKT W=1.62u L=40.00n
XX0 net053 A2 VDD VNW PHVT11LL_CKT W=1.62u L=40.00n
XX28 net053 A1 VDD VNW PHVT11LL_CKT W=1.62u L=40.00n
XX5 Z net053 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS AND3V8RD_12TH40
.SUBCKT AND3V8_12TH40 A1 A2 A3 Z VDD VSS
XX6 Z net053 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX2 net053 A1 net17 VPW NHVT11LL_CKT W=2.16u L=40.00n
XX9 net17 A2 net21 VPW NHVT11LL_CKT W=2.16u L=40.00n
XX8 net21 A3 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX1 net053 A3 VDD VNW PHVT11LL_CKT W=1.3u L=40.00n
XX0 net053 A2 VDD VNW PHVT11LL_CKT W=1.3u L=40.00n
XX28 net053 A1 VDD VNW PHVT11LL_CKT W=1.3u L=40.00n
XX5 Z net053 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS AND3V8_12TH40
.SUBCKT AND4V0_12TH40 A1 A2 A3 A4 Z VDD VSS
XX6 Z net032 VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX4 net032 A1 net26 VPW NHVT11LL_CKT W=310.00n L=40.00n
XX3 net26 A2 net30 VPW NHVT11LL_CKT W=310.00n L=40.00n
XX9 net30 A3 net34 VPW NHVT11LL_CKT W=310.00n L=40.00n
XX8 net34 A4 VSS VPW NHVT11LL_CKT W=310.00n L=40.00n
XX5 Z net032 VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
XX2 net032 A3 VDD VNW PHVT11LL_CKT W=150.00n L=40.00n
XX1 net032 A4 VDD VNW PHVT11LL_CKT W=150.00n L=40.00n
XX0 net032 A2 VDD VNW PHVT11LL_CKT W=150.00n L=40.00n
XX28 net032 A1 VDD VNW PHVT11LL_CKT W=150.00n L=40.00n
.ENDS AND4V0_12TH40
.SUBCKT AND4V10RD_12TH40 A1 A2 A3 A4 Z VDD VSS
XX6 Z net032 VSS VPW NHVT11LL_CKT W=2.7u L=40.00n
XX4 net032 A1 net26 VPW NHVT11LL_CKT W=6.1u L=40.00n
XX3 net26 A2 net30 VPW NHVT11LL_CKT W=6.1u L=40.00n
XX9 net30 A3 net34 VPW NHVT11LL_CKT W=6.1u L=40.00n
XX8 net34 A4 VSS VPW NHVT11LL_CKT W=6.1u L=40.00n
XX5 Z net032 VDD VNW PHVT11LL_CKT W=3.05u L=40.00n
XX2 net032 A3 VDD VNW PHVT11LL_CKT W=2.00u L=40.00n
XX1 net032 A4 VDD VNW PHVT11LL_CKT W=2.00u L=40.00n
XX0 net032 A2 VDD VNW PHVT11LL_CKT W=2.00u L=40.00n
XX28 net032 A1 VDD VNW PHVT11LL_CKT W=2.00u L=40.00n
.ENDS AND4V10RD_12TH40
.SUBCKT AND4V12_12TH40 A1 A2 A3 A4 Z VDD VSS
XX6 Z net032 VSS VPW NHVT11LL_CKT W=3.24u L=40.00n
XX4 net032 A1 net26 VPW NHVT11LL_CKT W=3.66u L=40.00n
XX3 net26 A2 net30 VPW NHVT11LL_CKT W=3.66u L=40.00n
XX9 net30 A3 net34 VPW NHVT11LL_CKT W=3.66u L=40.00n
XX8 net34 A4 VSS VPW NHVT11LL_CKT W=3.66u L=40.00n
XX5 Z net032 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX2 net032 A3 VDD VNW PHVT11LL_CKT W=1.8u L=40.00n
XX1 net032 A4 VDD VNW PHVT11LL_CKT W=1.8u L=40.00n
XX0 net032 A2 VDD VNW PHVT11LL_CKT W=1.8u L=40.00n
XX28 net032 A1 VDD VNW PHVT11LL_CKT W=1.8u L=40.00n
.ENDS AND4V12_12TH40
.SUBCKT AND4V16_12TH40 A1 A2 A3 A4 Z VDD VSS
XX6 Z net032 VSS VPW NHVT11LL_CKT W=4.32u L=40.00n
XX4 net032 A1 net26 VPW NHVT11LL_CKT W=4.88u L=40.00n
XX3 net26 A2 net30 VPW NHVT11LL_CKT W=4.88u L=40.00n
XX9 net30 A3 net34 VPW NHVT11LL_CKT W=4.88u L=40.00n
XX8 net34 A4 VSS VPW NHVT11LL_CKT W=4.88u L=40.00n
XX5 Z net032 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX2 net032 A3 VDD VNW PHVT11LL_CKT W=2.4u L=40.00n
XX1 net032 A4 VDD VNW PHVT11LL_CKT W=2.4u L=40.00n
XX0 net032 A2 VDD VNW PHVT11LL_CKT W=2.4u L=40.00n
XX28 net032 A1 VDD VNW PHVT11LL_CKT W=2.4u L=40.00n
.ENDS AND4V16_12TH40
.SUBCKT AND4V1RD_12TH40 A1 A2 A3 A4 Z VDD VSS
XX6 Z net032 VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX4 net032 A1 net26 VPW NHVT11LL_CKT W=850.00n L=40.00n
XX3 net26 A2 net30 VPW NHVT11LL_CKT W=850.00n L=40.00n
XX9 net30 A3 net34 VPW NHVT11LL_CKT W=850.00n L=40.00n
XX8 net34 A4 VSS VPW NHVT11LL_CKT W=850.00n L=40.00n
XX5 Z net032 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX2 net032 A3 VDD VNW PHVT11LL_CKT W=280.00n L=40.00n
XX1 net032 A4 VDD VNW PHVT11LL_CKT W=280.00n L=40.00n
XX0 net032 A2 VDD VNW PHVT11LL_CKT W=280.00n L=40.00n
XX28 net032 A1 VDD VNW PHVT11LL_CKT W=280.00n L=40.00n
.ENDS AND4V1RD_12TH40
.SUBCKT AND4V1_12TH40 A1 A2 A3 A4 Z VDD VSS
XX6 Z net032 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX4 net032 A1 net26 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX3 net26 A2 net30 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX9 net30 A3 net34 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX8 net34 A4 VSS VPW NHVT11LL_CKT W=430.00n L=40.00n
XX5 Z net032 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX2 net032 A3 VDD VNW PHVT11LL_CKT W=210.00n L=40.00n
XX1 net032 A4 VDD VNW PHVT11LL_CKT W=210.00n L=40.00n
XX0 net032 A2 VDD VNW PHVT11LL_CKT W=210.00n L=40.00n
XX28 net032 A1 VDD VNW PHVT11LL_CKT W=210.00n L=40.00n
.ENDS AND4V1_12TH40
.SUBCKT AND4V2RD_12TH40 A1 A2 A3 A4 Z VDD VSS
XX6 Z net032 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX4 net032 A1 net26 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX3 net26 A2 net30 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX9 net30 A3 net34 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX8 net34 A4 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX5 Z net032 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX2 net032 A3 VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX1 net032 A4 VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX0 net032 A2 VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX28 net032 A1 VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
.ENDS AND4V2RD_12TH40
.SUBCKT AND4V2_12TH40 A1 A2 A3 A4 Z VDD VSS
XX6 Z net032 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX4 net032 A1 net26 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX3 net26 A2 net30 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX9 net30 A3 net34 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX8 net34 A4 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX5 Z net032 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX2 net032 A3 VDD VNW PHVT11LL_CKT W=300.00n L=40.00n
XX1 net032 A4 VDD VNW PHVT11LL_CKT W=300.00n L=40.00n
XX0 net032 A2 VDD VNW PHVT11LL_CKT W=300.00n L=40.00n
XX28 net032 A1 VDD VNW PHVT11LL_CKT W=300.00n L=40.00n
.ENDS AND4V2_12TH40
.SUBCKT AND4V3_12TH40 A1 A2 A3 A4 Z VDD VSS
XX6 Z net032 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX4 net032 A1 net26 VPW NHVT11LL_CKT W=860.00n L=40.00n
XX3 net26 A2 net30 VPW NHVT11LL_CKT W=860.00n L=40.00n
XX9 net30 A3 net34 VPW NHVT11LL_CKT W=860.00n L=40.00n
XX8 net34 A4 VSS VPW NHVT11LL_CKT W=860.00n L=40.00n
XX5 Z net032 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX2 net032 A3 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX1 net032 A4 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX0 net032 A2 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX28 net032 A1 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
.ENDS AND4V3_12TH40
.SUBCKT AND4V4RD_12TH40 A1 A2 A3 A4 Z VDD VSS
XX6 Z net032 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX4 net032 A1 net26 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX3 net26 A2 net30 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX9 net30 A3 net34 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX8 net34 A4 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX5 Z net032 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX2 net032 A3 VDD VNW PHVT11LL_CKT W=800.00n L=40.00n
XX1 net032 A4 VDD VNW PHVT11LL_CKT W=800.00n L=40.00n
XX0 net032 A2 VDD VNW PHVT11LL_CKT W=800.00n L=40.00n
XX28 net032 A1 VDD VNW PHVT11LL_CKT W=800.00n L=40.00n
.ENDS AND4V4RD_12TH40
.SUBCKT AND4V4_12TH40 A1 A2 A3 A4 Z VDD VSS
XX6 Z net032 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX4 net032 A1 net26 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX3 net26 A2 net30 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX9 net30 A3 net34 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX8 net34 A4 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX5 Z net032 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX2 net032 A3 VDD VNW PHVT11LL_CKT W=600.00n L=40.00n
XX1 net032 A4 VDD VNW PHVT11LL_CKT W=600.00n L=40.00n
XX0 net032 A2 VDD VNW PHVT11LL_CKT W=600.00n L=40.00n
XX28 net032 A1 VDD VNW PHVT11LL_CKT W=600.00n L=40.00n
.ENDS AND4V4_12TH40
.SUBCKT AND4V6RD_12TH40 A1 A2 A3 A4 Z VDD VSS
XX6 Z net032 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX4 net032 A1 net26 VPW NHVT11LL_CKT W=3.66u L=40.00n
XX3 net26 A2 net30 VPW NHVT11LL_CKT W=3.66u L=40.00n
XX9 net30 A3 net34 VPW NHVT11LL_CKT W=3.66u L=40.00n
XX8 net34 A4 VSS VPW NHVT11LL_CKT W=3.66u L=40.00n
XX5 Z net032 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX2 net032 A3 VDD VNW PHVT11LL_CKT W=1.2u L=40.00n
XX1 net032 A4 VDD VNW PHVT11LL_CKT W=1.2u L=40.00n
XX0 net032 A2 VDD VNW PHVT11LL_CKT W=1.2u L=40.00n
XX28 net032 A1 VDD VNW PHVT11LL_CKT W=1.2u L=40.00n
.ENDS AND4V6RD_12TH40
.SUBCKT AND4V6_12TH40 A1 A2 A3 A4 Z VDD VSS
XX6 Z net032 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX4 net032 A1 net26 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX3 net26 A2 net30 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX9 net30 A3 net34 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX8 net34 A4 VSS VPW NHVT11LL_CKT W=1.83u L=40.00n
XX5 Z net032 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX2 net032 A3 VDD VNW PHVT11LL_CKT W=900.00n L=40.00n
XX1 net032 A4 VDD VNW PHVT11LL_CKT W=900.00n L=40.00n
XX0 net032 A2 VDD VNW PHVT11LL_CKT W=900.00n L=40.00n
XX28 net032 A1 VDD VNW PHVT11LL_CKT W=900.00n L=40.00n
.ENDS AND4V6_12TH40
.SUBCKT AND4V8RD_12TH40 A1 A2 A3 A4 Z VDD VSS
XX6 Z net032 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX4 net032 A1 net26 VPW NHVT11LL_CKT W=4.88u L=40.00n
XX3 net26 A2 net30 VPW NHVT11LL_CKT W=4.88u L=40.00n
XX9 net30 A3 net34 VPW NHVT11LL_CKT W=4.88u L=40.00n
XX8 net34 A4 VSS VPW NHVT11LL_CKT W=4.88u L=40.00n
XX5 Z net032 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX2 net032 A3 VDD VNW PHVT11LL_CKT W=1.6u L=40.00n
XX1 net032 A4 VDD VNW PHVT11LL_CKT W=1.6u L=40.00n
XX0 net032 A2 VDD VNW PHVT11LL_CKT W=1.6u L=40.00n
XX28 net032 A1 VDD VNW PHVT11LL_CKT W=1.6u L=40.00n
.ENDS AND4V8RD_12TH40
.SUBCKT AND4V8_12TH40 A1 A2 A3 A4 Z VDD VSS
XX6 Z net032 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX4 net032 A1 net26 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX3 net26 A2 net30 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX9 net30 A3 net34 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX8 net34 A4 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX5 Z net032 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX2 net032 A3 VDD VNW PHVT11LL_CKT W=1.2u L=40.00n
XX1 net032 A4 VDD VNW PHVT11LL_CKT W=1.2u L=40.00n
XX0 net032 A2 VDD VNW PHVT11LL_CKT W=1.2u L=40.00n
XX28 net032 A1 VDD VNW PHVT11LL_CKT W=1.2u L=40.00n
.ENDS AND4V8_12TH40
.SUBCKT AO1B2V0_12TH40 A1 A2 B Z VDD VSS
XX4 net29 B VSS VPW NHVT11LL_CKT W=0.305u L=40.00n
XX3 Z net9 net29 VPW NHVT11LL_CKT W=0.305u L=40.00n
XX9 net9 A1 net25 VPW NHVT11LL_CKT W=0.195u L=40.00n
XX8 net25 A2 VSS VPW NHVT11LL_CKT W=0.195u L=40.00n
XX2 Z net9 VDD VNW PHVT11LL_CKT W=0.295u L=40.00n
XX1 Z B VDD VNW PHVT11LL_CKT W=0.295u L=40.00n
XX0 net9 A1 VDD VNW PHVT11LL_CKT W=0.19u L=40.00n
XX28 net9 A2 VDD VNW PHVT11LL_CKT W=0.19u L=40.00n
.ENDS AO1B2V0_12TH40
.SUBCKT AO1B2V12_12TH40 A1 A2 B Z VDD VSS
XX4 net29 B VSS VPW NHVT11LL_CKT W=3.66u L=40.00n
XX3 Z net9 net29 VPW NHVT11LL_CKT W=3.66u L=40.00n
XX9 net9 A1 net25 VPW NHVT11LL_CKT W=1.695u L=40.00n
XX8 net25 A2 VSS VPW NHVT11LL_CKT W=1.695u L=40.00n
XX2 Z net9 VDD VNW PHVT11LL_CKT W=3.54u L=40.00n
XX1 Z B VDD VNW PHVT11LL_CKT W=3.54u L=40.00n
XX0 net9 A1 VDD VNW PHVT11LL_CKT W=1.635u L=40.00n
XX28 net9 A2 VDD VNW PHVT11LL_CKT W=1.635u L=40.00n
.ENDS AO1B2V12_12TH40
.SUBCKT AO1B2V1_12TH40 A1 A2 B Z VDD VSS
XX4 net29 B VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX3 Z net9 net29 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX9 net9 A1 net25 VPW NHVT11LL_CKT W=0.245u L=40.00n
XX8 net25 A2 VSS VPW NHVT11LL_CKT W=0.245u L=40.00n
XX2 Z net9 VDD VNW PHVT11LL_CKT W=0.415u L=40.00n
XX1 Z B VDD VNW PHVT11LL_CKT W=0.415u L=40.00n
XX0 net9 A1 VDD VNW PHVT11LL_CKT W=0.235u L=40.00n
XX28 net9 A2 VDD VNW PHVT11LL_CKT W=0.235u L=40.00n
.ENDS AO1B2V1_12TH40
.SUBCKT AO1B2V2_12TH40 A1 A2 B Z VDD VSS
XX4 net29 B VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX3 Z net9 net29 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX9 net9 A1 net25 VPW NHVT11LL_CKT W=315.00n L=40.00n
XX8 net25 A2 VSS VPW NHVT11LL_CKT W=315.00n L=40.00n
XX2 Z net9 VDD VNW PHVT11LL_CKT W=590.00n L=40.00n
XX1 Z B VDD VNW PHVT11LL_CKT W=590.00n L=40.00n
XX0 net9 A1 VDD VNW PHVT11LL_CKT W=305.00n L=40.00n
XX28 net9 A2 VDD VNW PHVT11LL_CKT W=305.00n L=40.00n
.ENDS AO1B2V2_12TH40
.SUBCKT AO1B2V3_12TH40 A1 A2 B Z VDD VSS
XX4 net29 B VSS VPW NHVT11LL_CKT W=0.86u L=40.00n
XX3 Z net9 net29 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX9 net9 A1 net25 VPW NHVT11LL_CKT W=0.42u L=40.00n
XX8 net25 A2 VSS VPW NHVT11LL_CKT W=0.42u L=40.00n
XX2 Z net9 VDD VNW PHVT11LL_CKT W=0.83u L=40.00n
XX1 Z B VDD VNW PHVT11LL_CKT W=0.83u L=40.00n
XX0 net9 A1 VDD VNW PHVT11LL_CKT W=0.41u L=40.00n
XX28 net9 A2 VDD VNW PHVT11LL_CKT W=0.41u L=40.00n
.ENDS AO1B2V3_12TH40
.SUBCKT AO1B2V4_12TH40 A1 A2 B Z VDD VSS
XX4 net29 B VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX3 Z net9 net29 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX9 net9 A1 net25 VPW NHVT11LL_CKT W=0.565u L=40.00n
XX8 net25 A2 VSS VPW NHVT11LL_CKT W=0.565u L=40.00n
XX2 Z net9 VDD VNW PHVT11LL_CKT W=1.18u L=40.00n
XX1 Z B VDD VNW PHVT11LL_CKT W=1.18u L=40.00n
XX0 net9 A1 VDD VNW PHVT11LL_CKT W=0.545u L=40.00n
XX28 net9 A2 VDD VNW PHVT11LL_CKT W=0.545u L=40.00n
.ENDS AO1B2V4_12TH40
.SUBCKT AO1B2V6_12TH40 A1 A2 B Z VDD VSS
XX4 net29 B VSS VPW NHVT11LL_CKT W=1.83u L=40.00n
XX3 Z net9 net29 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX9 net9 A1 net25 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX8 net25 A2 VSS VPW NHVT11LL_CKT W=0.86u L=40.00n
XX2 Z net9 VDD VNW PHVT11LL_CKT W=1.77u L=40.00n
XX1 Z B VDD VNW PHVT11LL_CKT W=1.77u L=40.00n
XX0 net9 A1 VDD VNW PHVT11LL_CKT W=0.83u L=40.00n
XX28 net9 A2 VDD VNW PHVT11LL_CKT W=0.83u L=40.00n
.ENDS AO1B2V6_12TH40
.SUBCKT AO1B2V8_12TH40 A1 A2 B Z VDD VSS
XX4 net29 B VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX3 Z net9 net29 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX9 net9 A1 net25 VPW NHVT11LL_CKT W=1.12u L=40.00n
XX8 net25 A2 VSS VPW NHVT11LL_CKT W=1.12u L=40.00n
XX2 Z net9 VDD VNW PHVT11LL_CKT W=2.36u L=40.00n
XX1 Z B VDD VNW PHVT11LL_CKT W=2.36u L=40.00n
XX0 net9 A1 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX28 net9 A2 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
.ENDS AO1B2V8_12TH40
.SUBCKT AO211V1_12TH40 A1 A2 B C Z VDD VSS
XX4 net028 C VSS VPW NHVT11LL_CKT W=150.00n L=40.00n
XX3 net028 B VSS VPW NHVT11LL_CKT W=150.00n L=40.00n
XX9 net028 A1 net18 VPW NHVT11LL_CKT W=270.00n L=40.00n
XX8 net18 A2 VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX5 Z net028 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX6 Z net028 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX2 net028 C net25 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX1 net25 B net34 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX0 net34 A2 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX28 net34 A1 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
.ENDS AO211V1_12TH40
.SUBCKT AO211V2_12TH40 A1 A2 B C Z VDD VSS
XX4 net028 C VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX3 net028 B VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX9 net028 A1 net18 VPW NHVT11LL_CKT W=380.00n L=40.00n
XX8 net18 A2 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX5 Z net028 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX6 Z net028 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX2 net028 C net25 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 net25 B net34 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX0 net34 A2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX28 net34 A1 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS AO211V2_12TH40
.SUBCKT AO211V4_12TH40 A1 A2 B C Z VDD VSS
XX4 net028 C VSS VPW NHVT11LL_CKT W=440.00n L=40.00n
XX3 net028 B VSS VPW NHVT11LL_CKT W=440.00n L=40.00n
XX9 net028 A1 net18 VPW NHVT11LL_CKT W=760.00n L=40.00n
XX8 net18 A2 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX5 Z net028 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX6 Z net028 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX2 net028 C net25 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 net25 B net34 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 net34 A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX28 net34 A1 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS AO211V4_12TH40
.SUBCKT AO211V8_12TH40 A1 A2 B C Z VDD VSS
XX4 net028 C VSS VPW NHVT11LL_CKT W=880.00n L=40.00n
XX3 net028 B VSS VPW NHVT11LL_CKT W=880.00n L=40.00n
XX9 net028 A1 net18 VPW NHVT11LL_CKT W=1.52u L=40.00n
XX8 net18 A2 VSS VPW NHVT11LL_CKT W=1.52u L=40.00n
XX5 Z net028 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX6 Z net028 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX2 net028 C net25 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 net25 B net34 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX0 net34 A2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX28 net34 A1 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS AO211V8_12TH40
.SUBCKT AO21BV0_12TH40 A1 A2 B Z VDD VSS
XX8 net5 A2 VSS VPW NHVT11LL_CKT W=0.195u L=40.00n
XX9 net071 A1 net5 VPW NHVT11LL_CKT W=0.195u L=40.00n
XX3 Z B net17 VPW NHVT11LL_CKT W=0.305u L=40.00n
XX4 net17 net071 VSS VPW NHVT11LL_CKT W=0.305u L=40.00n
XX28 net071 A2 VDD VNW PHVT11LL_CKT W=0.19u L=40.00n
XX0 net071 A1 VDD VNW PHVT11LL_CKT W=0.19u L=40.00n
XX1 Z B VDD VNW PHVT11LL_CKT W=0.295u L=40.00n
XX2 Z net071 VDD VNW PHVT11LL_CKT W=0.295u L=40.00n
.ENDS AO21BV0_12TH40
.SUBCKT AO21BV12_12TH40 A1 A2 B Z VDD VSS
XX8 net5 A2 VSS VPW NHVT11LL_CKT W=1.695u L=40.00n
XX9 net071 A1 net5 VPW NHVT11LL_CKT W=1.695u L=40.00n
XX3 Z B net17 VPW NHVT11LL_CKT W=3.66u L=40.00n
XX4 net17 net071 VSS VPW NHVT11LL_CKT W=3.66u L=40.00n
XX28 net071 A2 VDD VNW PHVT11LL_CKT W=1.635u L=40.00n
XX0 net071 A1 VDD VNW PHVT11LL_CKT W=1.635u L=40.00n
XX1 Z B VDD VNW PHVT11LL_CKT W=3.54u L=40.00n
XX2 Z net071 VDD VNW PHVT11LL_CKT W=3.54u L=40.00n
.ENDS AO21BV12_12TH40
.SUBCKT AO21BV1_12TH40 A1 A2 B Z VDD VSS
XX8 net5 A2 VSS VPW NHVT11LL_CKT W=0.245u L=40.00n
XX9 net071 A1 net5 VPW NHVT11LL_CKT W=0.245u L=40.00n
XX3 Z B net17 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX4 net17 net071 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX28 net071 A2 VDD VNW PHVT11LL_CKT W=0.235u L=40.00n
XX0 net071 A1 VDD VNW PHVT11LL_CKT W=0.235u L=40.00n
XX1 Z B VDD VNW PHVT11LL_CKT W=0.415u L=40.00n
XX2 Z net071 VDD VNW PHVT11LL_CKT W=0.415u L=40.00n
.ENDS AO21BV1_12TH40
.SUBCKT AO21BV2_12TH40 A1 A2 B Z VDD VSS
XX8 net5 A2 VSS VPW NHVT11LL_CKT W=315.00n L=40.00n
XX9 net071 A1 net5 VPW NHVT11LL_CKT W=315.00n L=40.00n
XX3 Z B net17 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX4 net17 net071 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX28 net071 A2 VDD VNW PHVT11LL_CKT W=305.00n L=40.00n
XX0 net071 A1 VDD VNW PHVT11LL_CKT W=305.00n L=40.00n
XX1 Z B VDD VNW PHVT11LL_CKT W=590.00n L=40.00n
XX2 Z net071 VDD VNW PHVT11LL_CKT W=590.00n L=40.00n
.ENDS AO21BV2_12TH40
.SUBCKT AO21BV3_12TH40 A1 A2 B Z VDD VSS
XX8 net5 A2 VSS VPW NHVT11LL_CKT W=0.42u L=40.00n
XX9 net071 A1 net5 VPW NHVT11LL_CKT W=0.42u L=40.00n
XX3 Z B net17 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX4 net17 net071 VSS VPW NHVT11LL_CKT W=0.86u L=40.00n
XX28 net071 A2 VDD VNW PHVT11LL_CKT W=0.41u L=40.00n
XX0 net071 A1 VDD VNW PHVT11LL_CKT W=0.41u L=40.00n
XX1 Z B VDD VNW PHVT11LL_CKT W=0.83u L=40.00n
XX2 Z net071 VDD VNW PHVT11LL_CKT W=0.83u L=40.00n
.ENDS AO21BV3_12TH40
.SUBCKT AO21BV4_12TH40 A1 A2 B Z VDD VSS
XX8 net5 A2 VSS VPW NHVT11LL_CKT W=0.565u L=40.00n
XX9 net071 A1 net5 VPW NHVT11LL_CKT W=0.565u L=40.00n
XX3 Z B net17 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX4 net17 net071 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX28 net071 A2 VDD VNW PHVT11LL_CKT W=0.545u L=40.00n
XX0 net071 A1 VDD VNW PHVT11LL_CKT W=0.545u L=40.00n
XX1 Z B VDD VNW PHVT11LL_CKT W=1.18u L=40.00n
XX2 Z net071 VDD VNW PHVT11LL_CKT W=1.18u L=40.00n
.ENDS AO21BV4_12TH40
.SUBCKT AO21BV6_12TH40 A1 A2 B Z VDD VSS
XX8 net5 A2 VSS VPW NHVT11LL_CKT W=0.86u L=40.00n
XX9 net071 A1 net5 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX3 Z B net17 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX4 net17 net071 VSS VPW NHVT11LL_CKT W=1.83u L=40.00n
XX28 net071 A2 VDD VNW PHVT11LL_CKT W=0.83u L=40.00n
XX0 net071 A1 VDD VNW PHVT11LL_CKT W=0.83u L=40.00n
XX1 Z B VDD VNW PHVT11LL_CKT W=1.77u L=40.00n
XX2 Z net071 VDD VNW PHVT11LL_CKT W=1.77u L=40.00n
.ENDS AO21BV6_12TH40
.SUBCKT AO21BV8_12TH40 A1 A2 B Z VDD VSS
XX8 net5 A2 VSS VPW NHVT11LL_CKT W=1.12u L=40.00n
XX9 net071 A1 net5 VPW NHVT11LL_CKT W=1.12u L=40.00n
XX3 Z B net17 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX4 net17 net071 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX28 net071 A2 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX0 net071 A1 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX1 Z B VDD VNW PHVT11LL_CKT W=2.36u L=40.00n
XX2 Z net071 VDD VNW PHVT11LL_CKT W=2.36u L=40.00n
.ENDS AO21BV8_12TH40
.SUBCKT AO21V0_12TH40 A1 A2 B Z VDD VSS
XX4 Z net048 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX2 net048 B VSS VPW NHVT11LL_CKT W=0.17u L=40.00n
XX9 net048 A1 net13 VPW NHVT11LL_CKT W=0.295u L=40.00n
XX8 net13 A2 VSS VPW NHVT11LL_CKT W=0.295u L=40.00n
XX3 Z net048 VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX1 net048 B net25 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX0 net25 A2 VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX28 net25 A1 VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
.ENDS AO21V0_12TH40
.SUBCKT AO21V12_12TH40 A1 A2 B Z VDD VSS
XX4 Z net048 VSS VPW NHVT11LL_CKT W=3.24u L=40.00n
XX2 net048 B VSS VPW NHVT11LL_CKT W=1.425u L=40.00n
XX9 net048 A1 net13 VPW NHVT11LL_CKT W=2.525u L=40.00n
XX8 net13 A2 VSS VPW NHVT11LL_CKT W=2.525u L=40.00n
XX3 Z net048 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX1 net048 B net25 VNW PHVT11LL_CKT W=3.05u L=40.00n
XX0 net25 A2 VDD VNW PHVT11LL_CKT W=3.05u L=40.00n
XX28 net25 A1 VDD VNW PHVT11LL_CKT W=3.05u L=40.00n
.ENDS AO21V12_12TH40
.SUBCKT AO21V1_12TH40 A1 A2 B Z VDD VSS
XX4 Z net048 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX2 net048 B VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX9 net048 A1 net13 VPW NHVT11LL_CKT W=0.365u L=40.00n
XX8 net13 A2 VSS VPW NHVT11LL_CKT W=0.365u L=40.00n
XX3 Z net048 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX1 net048 B net25 VNW PHVT11LL_CKT W=0.44u L=40.00n
XX0 net25 A2 VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX28 net25 A1 VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
.ENDS AO21V1_12TH40
.SUBCKT AO21V2_12TH40 A1 A2 B Z VDD VSS
XX4 Z net048 VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX2 net048 B VSS VPW NHVT11LL_CKT W=265.00n L=40.00n
XX9 net048 A1 net13 VPW NHVT11LL_CKT W=465.00n L=40.00n
XX8 net13 A2 VSS VPW NHVT11LL_CKT W=465.00n L=40.00n
XX3 Z net048 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 net048 B net25 VNW PHVT11LL_CKT W=565.00n L=40.00n
XX0 net25 A2 VDD VNW PHVT11LL_CKT W=565.00n L=40.00n
XX28 net25 A1 VDD VNW PHVT11LL_CKT W=565.00n L=40.00n
.ENDS AO21V2_12TH40
.SUBCKT AO21V3_12TH40 A1 A2 B Z VDD VSS
XX4 Z net048 VSS VPW NHVT11LL_CKT W=0.76u L=40.00n
XX2 net048 B VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX9 net048 A1 net13 VPW NHVT11LL_CKT W=0.67u L=40.00n
XX8 net13 A2 VSS VPW NHVT11LL_CKT W=0.67u L=40.00n
XX3 Z net048 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX1 net048 B net25 VNW PHVT11LL_CKT W=0.81u L=40.00n
XX0 net25 A2 VDD VNW PHVT11LL_CKT W=0.81u L=40.00n
XX28 net25 A1 VDD VNW PHVT11LL_CKT W=0.81u L=40.00n
.ENDS AO21V3_12TH40
.SUBCKT AO21V4_12TH40 A1 A2 B Z VDD VSS
XX4 Z net048 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX2 net048 B VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX9 net048 A1 net13 VPW NHVT11LL_CKT W=0.87u L=40.00n
XX8 net13 A2 VSS VPW NHVT11LL_CKT W=0.87u L=40.00n
XX3 Z net048 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 net048 B net25 VNW PHVT11LL_CKT W=1.05u L=40.00n
XX0 net25 A2 VDD VNW PHVT11LL_CKT W=1.05u L=40.00n
XX28 net25 A1 VDD VNW PHVT11LL_CKT W=1.05u L=40.00n
.ENDS AO21V4_12TH40
.SUBCKT AO21V6_12TH40 A1 A2 B Z VDD VSS
XX4 Z net048 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX2 net048 B VSS VPW NHVT11LL_CKT W=0.75u L=40.00n
XX9 net048 A1 net13 VPW NHVT11LL_CKT W=1.305u L=40.00n
XX8 net13 A2 VSS VPW NHVT11LL_CKT W=1.305u L=40.00n
XX3 Z net048 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX1 net048 B net25 VNW PHVT11LL_CKT W=1.575u L=40.00n
XX0 net25 A2 VDD VNW PHVT11LL_CKT W=1.575u L=40.00n
XX28 net25 A1 VDD VNW PHVT11LL_CKT W=1.575u L=40.00n
.ENDS AO21V6_12TH40
.SUBCKT AO21V8_12TH40 A1 A2 B Z VDD VSS
XX4 Z net048 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX2 net048 B VSS VPW NHVT11LL_CKT W=0.96u L=40.00n
XX9 net048 A1 net13 VPW NHVT11LL_CKT W=1.7u L=40.00n
XX8 net13 A2 VSS VPW NHVT11LL_CKT W=1.7u L=40.00n
XX3 Z net048 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 net048 B net25 VNW PHVT11LL_CKT W=2.04u L=40.00n
XX0 net25 A2 VDD VNW PHVT11LL_CKT W=2.04u L=40.00n
XX28 net25 A1 VDD VNW PHVT11LL_CKT W=2.04u L=40.00n
.ENDS AO21V8_12TH40
.SUBCKT AO221V1_12TH40 A1 A2 B1 B2 C Z VDD VSS
XX4 net024 C VSS VPW NHVT11LL_CKT W=150.00n L=40.00n
XX2 net024 B1 net31 VPW NHVT11LL_CKT W=270.00n L=40.00n
XX9 net024 A1 net43 VPW NHVT11LL_CKT W=270.00n L=40.00n
XX8 net43 A2 VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX7 Z net024 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX3 net31 B2 VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX10 Z net024 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX6 net26 A1 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX5 net26 A2 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX1 net024 C net23 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX0 net23 B2 net26 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX28 net23 B1 net26 VNW PHVT11LL_CKT W=430.00n L=40.00n
.ENDS AO221V1_12TH40
.SUBCKT AO221V2_12TH40 A1 A2 B1 B2 C Z VDD VSS
XX4 net024 C VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX2 net024 B1 net31 VPW NHVT11LL_CKT W=380.00n L=40.00n
XX9 net024 A1 net43 VPW NHVT11LL_CKT W=380.00n L=40.00n
XX8 net43 A2 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX7 Z net024 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX3 net31 B2 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX10 Z net024 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX6 net26 A1 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX5 net26 A2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 net024 C net23 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX0 net23 B2 net26 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX28 net23 B1 net26 VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS AO221V2_12TH40
.SUBCKT AO221V4_12TH40 A1 A2 B1 B2 C Z VDD VSS
XX4 net024 C VSS VPW NHVT11LL_CKT W=440.00n L=40.00n
XX2 net024 B1 net31 VPW NHVT11LL_CKT W=760.00n L=40.00n
XX9 net024 A1 net43 VPW NHVT11LL_CKT W=760.00n L=40.00n
XX8 net43 A2 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX7 Z net024 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX3 net31 B2 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX10 Z net024 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX6 net26 A1 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX5 net26 A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 net024 C net23 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 net23 B2 net26 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX28 net23 B1 net26 VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS AO221V4_12TH40
.SUBCKT AO221V8_12TH40 A1 A2 B1 B2 C Z VDD VSS
XX4 net024 C VSS VPW NHVT11LL_CKT W=880.00n L=40.00n
XX2 net024 B1 net31 VPW NHVT11LL_CKT W=1.52u L=40.00n
XX9 net024 A1 net43 VPW NHVT11LL_CKT W=1.52u L=40.00n
XX8 net43 A2 VSS VPW NHVT11LL_CKT W=1.52u L=40.00n
XX7 Z net024 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX3 net31 B2 VSS VPW NHVT11LL_CKT W=1.52u L=40.00n
XX10 Z net024 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX6 net26 A1 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX5 net26 A2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 net024 C net23 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX0 net23 B2 net26 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX28 net23 B1 net26 VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS AO221V8_12TH40
.SUBCKT AO222V1_12TH40 A1 A2 B1 B2 C1 C2 Z VDD VSS
XX11 Z net049 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX7 net8 C2 VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX3 net12 B2 VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX8 net16 A2 VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX9 net049 A1 net16 VPW NHVT11LL_CKT W=270.00n L=40.00n
XX2 net049 B1 net12 VPW NHVT11LL_CKT W=270.00n L=40.00n
XX4 net049 C1 net8 VPW NHVT11LL_CKT W=270.00n L=40.00n
XX12 Z net049 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX10 net049 C2 net39 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX28 net39 B1 net43 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX0 net39 B2 net43 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX1 net049 C1 net39 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX5 net43 A2 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX6 net43 A1 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
.ENDS AO222V1_12TH40
.SUBCKT AO222V2_12TH40 A1 A2 B1 B2 C1 C2 Z VDD VSS
XX11 Z net049 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX7 net8 C2 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX3 net12 B2 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX8 net16 A2 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX9 net049 A1 net16 VPW NHVT11LL_CKT W=380.00n L=40.00n
XX2 net049 B1 net12 VPW NHVT11LL_CKT W=380.00n L=40.00n
XX4 net049 C1 net8 VPW NHVT11LL_CKT W=380.00n L=40.00n
XX12 Z net049 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX10 net049 C2 net39 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX28 net39 B1 net43 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX0 net39 B2 net43 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 net049 C1 net39 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX5 net43 A2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX6 net43 A1 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS AO222V2_12TH40
.SUBCKT AO222V4_12TH40 A1 A2 B1 B2 C1 C2 Z VDD VSS
XX11 Z net049 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX7 net8 C2 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX3 net12 B2 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX8 net16 A2 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX9 net049 A1 net16 VPW NHVT11LL_CKT W=760.00n L=40.00n
XX2 net049 B1 net12 VPW NHVT11LL_CKT W=760.00n L=40.00n
XX4 net049 C1 net8 VPW NHVT11LL_CKT W=760.00n L=40.00n
XX12 Z net049 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX10 net049 C2 net39 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX28 net39 B1 net43 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 net39 B2 net43 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 net049 C1 net39 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX5 net43 A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX6 net43 A1 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS AO222V4_12TH40
.SUBCKT AO222V8_12TH40 A1 A2 B1 B2 C1 C2 Z VDD VSS
XX11 Z net049 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX7 net8 C2 VSS VPW NHVT11LL_CKT W=1.52u L=40.00n
XX3 net12 B2 VSS VPW NHVT11LL_CKT W=1.52u L=40.00n
XX8 net16 A2 VSS VPW NHVT11LL_CKT W=1.52u L=40.00n
XX9 net049 A1 net16 VPW NHVT11LL_CKT W=1.52u L=40.00n
XX2 net049 B1 net12 VPW NHVT11LL_CKT W=1.52u L=40.00n
XX4 net049 C1 net8 VPW NHVT11LL_CKT W=1.52u L=40.00n
XX12 Z net049 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX10 net049 C2 net39 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX28 net39 B1 net43 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX0 net39 B2 net43 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 net049 C1 net39 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX5 net43 A2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX6 net43 A1 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS AO222V8_12TH40
.SUBCKT AO22V0_12TH40 A1 A2 B1 B2 Z VDD VSS
XX6 Z net068 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX4 net6 B2 VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX3 net068 B1 net6 VPW NHVT11LL_CKT W=0.31u L=40.00n
XX9 net068 A1 net18 VPW NHVT11LL_CKT W=0.31u L=40.00n
XX8 net18 A2 VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX5 Z net068 VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX2 net068 B2 net29 VNW PHVT11LL_CKT W=0.37u L=40.00n
XX1 net068 B1 net29 VNW PHVT11LL_CKT W=0.37u L=40.00n
XX0 net29 A2 VDD VNW PHVT11LL_CKT W=0.37u L=40.00n
XX28 net29 A1 VDD VNW PHVT11LL_CKT W=0.37u L=40.00n
.ENDS AO22V0_12TH40
.SUBCKT AO22V12_12TH40 A1 A2 B1 B2 Z VDD VSS
XX6 Z net068 VSS VPW NHVT11LL_CKT W=3.24u L=40.00n
XX4 net6 B2 VSS VPW NHVT11LL_CKT W=2.79u L=40.00n
XX3 net068 B1 net6 VPW NHVT11LL_CKT W=2.79u L=40.00n
XX9 net068 A1 net18 VPW NHVT11LL_CKT W=2.79u L=40.00n
XX8 net18 A2 VSS VPW NHVT11LL_CKT W=2.79u L=40.00n
XX5 Z net068 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX2 net068 B2 net29 VNW PHVT11LL_CKT W=3.36u L=40.00n
XX1 net068 B1 net29 VNW PHVT11LL_CKT W=3.36u L=40.00n
XX0 net29 A2 VDD VNW PHVT11LL_CKT W=3.36u L=40.00n
XX28 net29 A1 VDD VNW PHVT11LL_CKT W=3.36u L=40.00n
.ENDS AO22V12_12TH40
.SUBCKT AO22V1_12TH40 A1 A2 B1 B2 Z VDD VSS
XX6 Z net068 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX4 net6 B2 VSS VPW NHVT11LL_CKT W=0.375u L=40.00n
XX3 net068 B1 net6 VPW NHVT11LL_CKT W=0.375u L=40.00n
XX9 net068 A1 net18 VPW NHVT11LL_CKT W=0.375u L=40.00n
XX8 net18 A2 VSS VPW NHVT11LL_CKT W=0.375u L=40.00n
XX5 Z net068 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX2 net068 B2 net29 VNW PHVT11LL_CKT W=0.455u L=40.00n
XX1 net068 B1 net29 VNW PHVT11LL_CKT W=0.455u L=40.00n
XX0 net29 A2 VDD VNW PHVT11LL_CKT W=0.455u L=40.00n
XX28 net29 A1 VDD VNW PHVT11LL_CKT W=0.455u L=40.00n
.ENDS AO22V1_12TH40
.SUBCKT AO22V2_12TH40 A1 A2 B1 B2 Z VDD VSS
XX6 Z net068 VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX4 net6 B2 VSS VPW NHVT11LL_CKT W=480.00n L=40.00n
XX3 net068 B1 net6 VPW NHVT11LL_CKT W=480.00n L=40.00n
XX9 net068 A1 net18 VPW NHVT11LL_CKT W=480.00n L=40.00n
XX8 net18 A2 VSS VPW NHVT11LL_CKT W=480.00n L=40.00n
XX5 Z net068 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX2 net068 B2 net29 VNW PHVT11LL_CKT W=580.00n L=40.00n
XX1 net068 B1 net29 VNW PHVT11LL_CKT W=580.00n L=40.00n
XX0 net29 A2 VDD VNW PHVT11LL_CKT W=580.00n L=40.00n
XX28 net29 A1 VDD VNW PHVT11LL_CKT W=580.00n L=40.00n
.ENDS AO22V2_12TH40
.SUBCKT AO22V3_12TH40 A1 A2 B1 B2 Z VDD VSS
XX6 Z net068 VSS VPW NHVT11LL_CKT W=0.76u L=40.00n
XX4 net6 B2 VSS VPW NHVT11LL_CKT W=0.75u L=40.00n
XX3 net068 B1 net6 VPW NHVT11LL_CKT W=0.75u L=40.00n
XX9 net068 A1 net18 VPW NHVT11LL_CKT W=0.75u L=40.00n
XX8 net18 A2 VSS VPW NHVT11LL_CKT W=0.75u L=40.00n
XX5 Z net068 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX2 net068 B2 net29 VNW PHVT11LL_CKT W=0.9u L=40.00n
XX1 net068 B1 net29 VNW PHVT11LL_CKT W=0.9u L=40.00n
XX0 net29 A2 VDD VNW PHVT11LL_CKT W=0.9u L=40.00n
XX28 net29 A1 VDD VNW PHVT11LL_CKT W=0.9u L=40.00n
.ENDS AO22V3_12TH40
.SUBCKT AO22V4_12TH40 A1 A2 B1 B2 Z VDD VSS
XX6 Z net068 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX4 net6 B2 VSS VPW NHVT11LL_CKT W=0.95u L=40.00n
XX3 net068 B1 net6 VPW NHVT11LL_CKT W=0.95u L=40.00n
XX9 net068 A1 net18 VPW NHVT11LL_CKT W=0.95u L=40.00n
XX8 net18 A2 VSS VPW NHVT11LL_CKT W=0.95u L=40.00n
XX5 Z net068 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX2 net068 B2 net29 VNW PHVT11LL_CKT W=1.15u L=40.00n
XX1 net068 B1 net29 VNW PHVT11LL_CKT W=1.15u L=40.00n
XX0 net29 A2 VDD VNW PHVT11LL_CKT W=1.15u L=40.00n
XX28 net29 A1 VDD VNW PHVT11LL_CKT W=1.15u L=40.00n
.ENDS AO22V4_12TH40
.SUBCKT AO22V6_12TH40 A1 A2 B1 B2 Z VDD VSS
XX6 Z net068 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX4 net6 B2 VSS VPW NHVT11LL_CKT W=1.47u L=40.00n
XX3 net068 B1 net6 VPW NHVT11LL_CKT W=1.47u L=40.00n
XX9 net068 A1 net18 VPW NHVT11LL_CKT W=1.47u L=40.00n
XX8 net18 A2 VSS VPW NHVT11LL_CKT W=1.47u L=40.00n
XX5 Z net068 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX2 net068 B2 net29 VNW PHVT11LL_CKT W=1.77u L=40.00n
XX1 net068 B1 net29 VNW PHVT11LL_CKT W=1.77u L=40.00n
XX0 net29 A2 VDD VNW PHVT11LL_CKT W=1.77u L=40.00n
XX28 net29 A1 VDD VNW PHVT11LL_CKT W=1.77u L=40.00n
.ENDS AO22V6_12TH40
.SUBCKT AO22V8_12TH40 A1 A2 B1 B2 Z VDD VSS
XX6 Z net068 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX4 net6 B2 VSS VPW NHVT11LL_CKT W=1.88u L=40.00n
XX3 net068 B1 net6 VPW NHVT11LL_CKT W=1.88u L=40.00n
XX9 net068 A1 net18 VPW NHVT11LL_CKT W=1.88u L=40.00n
XX8 net18 A2 VSS VPW NHVT11LL_CKT W=1.88u L=40.00n
XX5 Z net068 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX2 net068 B2 net29 VNW PHVT11LL_CKT W=2.28u L=40.00n
XX1 net068 B1 net29 VNW PHVT11LL_CKT W=2.28u L=40.00n
XX0 net29 A2 VDD VNW PHVT11LL_CKT W=2.28u L=40.00n
XX28 net29 A1 VDD VNW PHVT11LL_CKT W=2.28u L=40.00n
.ENDS AO22V8_12TH40
.SUBCKT AO31V1_12TH40 A1 A2 A3 B Z VDD VSS
XX3 net22 A3 VSS VPW NHVT11LL_CKT W=430.00n L=40.00n
XX2 net026 B VSS VPW NHVT11LL_CKT W=190.00n L=40.00n
XX9 net026 A1 net34 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX8 net34 A2 net22 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX6 Z net026 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX5 Z net026 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX4 net6 A3 VDD VNW PHVT11LL_CKT W=380.00n L=40.00n
XX1 net026 B net6 VNW PHVT11LL_CKT W=380.00n L=40.00n
XX0 net6 A2 VDD VNW PHVT11LL_CKT W=380.00n L=40.00n
XX28 net6 A1 VDD VNW PHVT11LL_CKT W=380.00n L=40.00n
.ENDS AO31V1_12TH40
.SUBCKT AO31V2_12TH40 A1 A2 A3 B Z VDD VSS
XX3 net22 A3 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX2 net026 B VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX9 net026 A1 net34 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX8 net34 A2 net22 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX6 Z net026 VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX5 Z net026 VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX4 net6 A3 VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX1 net026 B net6 VNW PHVT11LL_CKT W=540.00n L=40.00n
XX0 net6 A2 VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX28 net6 A1 VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
.ENDS AO31V2_12TH40
.SUBCKT AO31V4_12TH40 A1 A2 A3 B Z VDD VSS
XX3 net22 A3 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX2 net026 B VSS VPW NHVT11LL_CKT W=1u L=40.00n
XX9 net026 A1 net34 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX8 net34 A2 net22 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX6 Z net026 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX5 Z net026 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX4 net6 A3 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX1 net026 B net6 VNW PHVT11LL_CKT W=1.08u L=40.00n
XX0 net6 A2 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX28 net6 A1 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
.ENDS AO31V4_12TH40
.SUBCKT AO31V8_12TH40 A1 A2 A3 B Z VDD VSS
XX3 net22 A3 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX2 net026 B VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX9 net026 A1 net34 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX8 net34 A2 net22 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX6 Z net026 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX5 Z net026 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX4 net6 A3 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
XX1 net026 B net6 VNW PHVT11LL_CKT W=2.16u L=40.00n
XX0 net6 A2 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
XX28 net6 A1 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
.ENDS AO31V8_12TH40
.SUBCKT AO32V1_12TH40 A1 A2 A3 B1 B2 Z VDD VSS
XX7 Z net035 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX5 net056 B2 VSS VPW NHVT11LL_CKT W=330.00n L=40.00n
XX8 net6 A2 net18 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX9 net035 A1 net6 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX2 net035 B1 net056 VPW NHVT11LL_CKT W=330.00n L=40.00n
XX3 net18 A3 VSS VPW NHVT11LL_CKT W=430.00n L=40.00n
XX10 Z net035 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX6 net035 B1 net34 VNW PHVT11LL_CKT W=380.00n L=40.00n
XX1 net035 B2 net34 VNW PHVT11LL_CKT W=380.00n L=40.00n
XX0 net34 A2 VDD VNW PHVT11LL_CKT W=380.00n L=40.00n
XX4 net34 A3 VDD VNW PHVT11LL_CKT W=380.00n L=40.00n
XX28 net34 A1 VDD VNW PHVT11LL_CKT W=380.00n L=40.00n
.ENDS AO32V1_12TH40
.SUBCKT AO32V2_12TH40 A1 A2 A3 B1 B2 Z VDD VSS
XX7 Z net035 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX5 net056 B2 VSS VPW NHVT11LL_CKT W=460.00n L=40.00n
XX8 net6 A2 net18 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX9 net035 A1 net6 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX2 net035 B1 net056 VPW NHVT11LL_CKT W=460.00n L=40.00n
XX3 net18 A3 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX10 Z net035 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX6 net035 B1 net34 VNW PHVT11LL_CKT W=540.00n L=40.00n
XX1 net035 B2 net34 VNW PHVT11LL_CKT W=540.00n L=40.00n
XX0 net34 A2 VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX4 net34 A3 VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX28 net34 A1 VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
.ENDS AO32V2_12TH40
.SUBCKT AO32V4_12TH40 A1 A2 A3 B1 B2 Z VDD VSS
XX7 Z net035 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX5 net056 B2 VSS VPW NHVT11LL_CKT W=920.00n L=40.00n
XX8 net6 A2 net18 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX9 net035 A1 net6 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX2 net035 B1 net056 VPW NHVT11LL_CKT W=920.00n L=40.00n
XX3 net18 A3 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX10 Z net035 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX6 net035 B1 net34 VNW PHVT11LL_CKT W=1.08u L=40.00n
XX1 net035 B2 net34 VNW PHVT11LL_CKT W=1.08u L=40.00n
XX0 net34 A2 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX4 net34 A3 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX28 net34 A1 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
.ENDS AO32V4_12TH40
.SUBCKT AO32V8_12TH40 A1 A2 A3 B1 B2 Z VDD VSS
XX7 Z net035 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX5 net056 B2 VSS VPW NHVT11LL_CKT W=1.84u L=40.00n
XX8 net6 A2 net18 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX9 net035 A1 net6 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX2 net035 B1 net056 VPW NHVT11LL_CKT W=1.84u L=40.00n
XX3 net18 A3 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX10 Z net035 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX6 net035 B1 net34 VNW PHVT11LL_CKT W=2.16u L=40.00n
XX1 net035 B2 net34 VNW PHVT11LL_CKT W=2.16u L=40.00n
XX0 net34 A2 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
XX4 net34 A3 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
XX28 net34 A1 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
.ENDS AO32V8_12TH40
.SUBCKT AO33V1_12TH40 A1 A2 A3 B1 B2 B3 Z VDD VSS
XX7 Z net035 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX11 net028 B3 VSS VPW NHVT11LL_CKT W=430.00n L=40.00n
XX5 net056 B2 net028 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX8 net6 A2 net18 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX9 net035 A1 net6 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX2 net035 B1 net056 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX3 net18 A3 VSS VPW NHVT11LL_CKT W=430.00n L=40.00n
XX10 Z net035 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX12 net035 B3 net34 VNW PHVT11LL_CKT W=380.00n L=40.00n
XX6 net035 B1 net34 VNW PHVT11LL_CKT W=380.00n L=40.00n
XX1 net035 B2 net34 VNW PHVT11LL_CKT W=380.00n L=40.00n
XX0 net34 A2 VDD VNW PHVT11LL_CKT W=380.00n L=40.00n
XX4 net34 A3 VDD VNW PHVT11LL_CKT W=380.00n L=40.00n
XX28 net34 A1 VDD VNW PHVT11LL_CKT W=380.00n L=40.00n
.ENDS AO33V1_12TH40
.SUBCKT AO33V2_12TH40 A1 A2 A3 B1 B2 B3 Z VDD VSS
XX0 net43 A2 VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX4 net43 A3 VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX28 net43 A1 VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX10 Z net40 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX12 net40 B3 net43 VNW PHVT11LL_CKT W=540.00n L=40.00n
XX6 net40 B1 net43 VNW PHVT11LL_CKT W=540.00n L=40.00n
XX1 net40 B2 net43 VNW PHVT11LL_CKT W=540.00n L=40.00n
XX7 Z net40 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX3 net52 A3 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX11 net72 B3 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX5 net68 B2 net72 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX8 net64 A2 net52 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX9 net40 A1 net64 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX2 net40 B1 net68 VPW NHVT11LL_CKT W=610.00n L=40.00n
.ENDS AO33V2_12TH40
.SUBCKT AO33V4_12TH40 A1 A2 A3 B1 B2 B3 Z VDD VSS
XX0 net43 A2 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX4 net43 A3 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX28 net43 A1 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX10 Z net40 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX12 net40 B3 net43 VNW PHVT11LL_CKT W=1.08u L=40.00n
XX6 net40 B1 net43 VNW PHVT11LL_CKT W=1.08u L=40.00n
XX1 net40 B2 net43 VNW PHVT11LL_CKT W=1.08u L=40.00n
XX7 Z net40 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX3 net52 A3 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX11 net72 B3 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX5 net68 B2 net72 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX8 net64 A2 net52 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX9 net40 A1 net64 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX2 net40 B1 net68 VPW NHVT11LL_CKT W=1.22u L=40.00n
.ENDS AO33V4_12TH40
.SUBCKT AO33V8_12TH40 A1 A2 A3 B1 B2 B3 Z VDD VSS
XX0 net43 A2 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
XX4 net43 A3 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
XX28 net43 A1 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
XX10 Z net40 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX12 net40 B3 net43 VNW PHVT11LL_CKT W=2.16u L=40.00n
XX6 net40 B1 net43 VNW PHVT11LL_CKT W=2.16u L=40.00n
XX1 net40 B2 net43 VNW PHVT11LL_CKT W=2.16u L=40.00n
XX7 Z net40 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX3 net52 A3 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX11 net72 B3 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX5 net68 B2 net72 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX8 net64 A2 net52 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX9 net40 A1 net64 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX2 net40 B1 net68 VPW NHVT11LL_CKT W=2.44u L=40.00n
.ENDS AO33V8_12TH40
.SUBCKT AOA211V1_12TH40 A1 A2 B C Z VDD VSS
XX7 Z net044 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX3 net044 C net30 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX2 net30 B VSS VPW NHVT11LL_CKT W=330.00n L=40.00n
XX9 net30 A1 net34 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX8 net34 A2 VSS VPW NHVT11LL_CKT W=430.00n L=40.00n
XX10 Z net044 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX4 net044 C VDD VNW PHVT11LL_CKT W=230.00n L=40.00n
XX1 net044 B net18 VNW PHVT11LL_CKT W=380.00n L=40.00n
XX0 net18 A1 VDD VNW PHVT11LL_CKT W=380.00n L=40.00n
XX28 net18 A2 VDD VNW PHVT11LL_CKT W=380.00n L=40.00n
.ENDS AOA211V1_12TH40
.SUBCKT AOA211V2_12TH40 A1 A2 B C Z VDD VSS
XX7 Z net044 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX3 net044 C net30 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX2 net30 B VSS VPW NHVT11LL_CKT W=460.00n L=40.00n
XX9 net30 A1 net34 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX8 net34 A2 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX10 Z net044 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX4 net044 C VDD VNW PHVT11LL_CKT W=0.32u L=40.00n
XX1 net044 B net18 VNW PHVT11LL_CKT W=540.00n L=40.00n
XX0 net18 A1 VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX28 net18 A2 VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
.ENDS AOA211V2_12TH40
.SUBCKT AOA211V4_12TH40 A1 A2 B C Z VDD VSS
XX7 Z net044 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX3 net044 C net30 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX2 net30 B VSS VPW NHVT11LL_CKT W=920.00n L=40.00n
XX9 net30 A1 net34 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX8 net34 A2 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX10 Z net044 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX4 net044 C VDD VNW PHVT11LL_CKT W=620.00n L=40.00n
XX1 net044 B net18 VNW PHVT11LL_CKT W=1.08u L=40.00n
XX0 net18 A1 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX28 net18 A2 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
.ENDS AOA211V4_12TH40
.SUBCKT AOA211V8_12TH40 A1 A2 B C Z VDD VSS
XX7 Z net044 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX3 net044 C net30 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX2 net30 B VSS VPW NHVT11LL_CKT W=1.84u L=40.00n
XX9 net30 A1 net34 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX8 net34 A2 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX10 Z net044 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX4 net044 C VDD VNW PHVT11LL_CKT W=1.24u L=40.00n
XX1 net044 B net18 VNW PHVT11LL_CKT W=2.16u L=40.00n
XX0 net18 A1 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
XX28 net18 A2 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
.ENDS AOA211V8_12TH40
.SUBCKT AOAI211V0_12TH40 A1 A2 B C ZN VDD VSS
XX3 ZN C net30 VPW NHVT11LL_CKT W=0.305u L=40.00n
XX2 net30 B VSS VPW NHVT11LL_CKT W=0.22u L=40.00n
XX9 net30 A1 net34 VPW NHVT11LL_CKT W=0.305u L=40.00n
XX8 net34 A2 VSS VPW NHVT11LL_CKT W=0.305u L=40.00n
XX4 ZN C VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX1 ZN B net18 VNW PHVT11LL_CKT W=0.27u L=40.00n
XX0 net18 A1 VDD VNW PHVT11LL_CKT W=0.27u L=40.00n
XX28 net18 A2 VDD VNW PHVT11LL_CKT W=0.27u L=40.00n
.ENDS AOAI211V0_12TH40
.SUBCKT AOAI211V12_12TH40 A1 A2 B C ZN VDD VSS
XX3 ZN C net30 VPW NHVT11LL_CKT W=3.66u L=40.00n
XX2 net30 B VSS VPW NHVT11LL_CKT W=2.64u L=40.00n
XX9 net30 A1 net34 VPW NHVT11LL_CKT W=3.66u L=40.00n
XX8 net34 A2 VSS VPW NHVT11LL_CKT W=3.66u L=40.00n
XX4 ZN C VDD VNW PHVT11LL_CKT W=1.71u L=40.00n
XX1 ZN B net18 VNW PHVT11LL_CKT W=3.24u L=40.00n
XX0 net18 A1 VDD VNW PHVT11LL_CKT W=3.24u L=40.00n
XX28 net18 A2 VDD VNW PHVT11LL_CKT W=3.24u L=40.00n
.ENDS AOAI211V12_12TH40
.SUBCKT AOAI211V1_12TH40 A1 A2 B C ZN VDD VSS
XX3 ZN C net30 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX2 net30 B VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX9 net30 A1 net34 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX8 net34 A2 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX4 ZN C VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX1 ZN B net18 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX0 net18 A1 VDD VNW PHVT11LL_CKT W=0.38u L=40.00n
XX28 net18 A2 VDD VNW PHVT11LL_CKT W=0.38u L=40.00n
.ENDS AOAI211V1_12TH40
.SUBCKT AOAI211V2_12TH40 A1 A2 B C ZN VDD VSS
XX3 ZN C net30 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX2 net30 B VSS VPW NHVT11LL_CKT W=440.00n L=40.00n
XX9 net30 A1 net34 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX8 net34 A2 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX4 ZN C VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX1 ZN B net18 VNW PHVT11LL_CKT W=0.54u L=40.00n
XX0 net18 A1 VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX28 net18 A2 VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
.ENDS AOAI211V2_12TH40
.SUBCKT AOAI211V3_12TH40 A1 A2 B C ZN VDD VSS
XX3 ZN C net30 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX2 net30 B VSS VPW NHVT11LL_CKT W=0.62u L=40.00n
XX9 net30 A1 net34 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX8 net34 A2 VSS VPW NHVT11LL_CKT W=0.86u L=40.00n
XX4 ZN C VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX1 ZN B net18 VNW PHVT11LL_CKT W=0.76u L=40.00n
XX0 net18 A1 VDD VNW PHVT11LL_CKT W=0.76u L=40.00n
XX28 net18 A2 VDD VNW PHVT11LL_CKT W=0.76u L=40.00n
.ENDS AOAI211V3_12TH40
.SUBCKT AOAI211V4_12TH40 A1 A2 B C ZN VDD VSS
XX3 ZN C net30 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX2 net30 B VSS VPW NHVT11LL_CKT W=0.88u L=40.00n
XX9 net30 A1 net34 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX8 net34 A2 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX4 ZN C VDD VNW PHVT11LL_CKT W=0.57u L=40.00n
XX1 ZN B net18 VNW PHVT11LL_CKT W=1.08u L=40.00n
XX0 net18 A1 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX28 net18 A2 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
.ENDS AOAI211V4_12TH40
.SUBCKT AOAI211V6_12TH40 A1 A2 B C ZN VDD VSS
XX3 ZN C net30 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX2 net30 B VSS VPW NHVT11LL_CKT W=1.32u L=40.00n
XX9 net30 A1 net34 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX8 net34 A2 VSS VPW NHVT11LL_CKT W=1.83u L=40.00n
XX4 ZN C VDD VNW PHVT11LL_CKT W=0.855u L=40.00n
XX1 ZN B net18 VNW PHVT11LL_CKT W=1.62u L=40.00n
XX0 net18 A1 VDD VNW PHVT11LL_CKT W=1.62u L=40.00n
XX28 net18 A2 VDD VNW PHVT11LL_CKT W=1.62u L=40.00n
.ENDS AOAI211V6_12TH40
.SUBCKT AOAI211V8_12TH40 A1 A2 B C ZN VDD VSS
XX3 ZN C net30 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX2 net30 B VSS VPW NHVT11LL_CKT W=1.76u L=40.00n
XX9 net30 A1 net34 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX8 net34 A2 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX4 ZN C VDD VNW PHVT11LL_CKT W=1.14u L=40.00n
XX1 ZN B net18 VNW PHVT11LL_CKT W=2.16u L=40.00n
XX0 net18 A1 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
XX28 net18 A2 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
.ENDS AOAI211V8_12TH40
.SUBCKT AOAOAOI211111V1_12TH40 A1 A2 B C D E F ZN VDD VSS
XX14 ZN E net_21 VPW NHVT11LL_CKT W=380.00n L=40.00n
XX13 ZN F VSS VPW NHVT11LL_CKT W=190.00n L=40.00n
XX12 net_21 D VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX10 net_21 C net_29 VPW NHVT11LL_CKT W=380.00n L=40.00n
XX9 net_29 B VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX8 net_29 A1 net4 VPW NHVT11LL_CKT W=380.00n L=40.00n
XX7 net4 A2 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX6 net_64 E VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
XX5 net_60 C VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX4 net3 A2 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX3 net3 A1 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX2 net_60 B net3 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX1 net_64 D net_60 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX0 ZN F net_64 VNW PHVT11LL_CKT W=430.00n L=40.00n
.ENDS AOAOAOI211111V1_12TH40
.SUBCKT AOAOAOI211111V2_12TH40 A1 A2 B C D E F ZN VDD VSS
XX6 net_71 E VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX5 net_75 C VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX4 net3 A2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX3 net3 A1 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX2 net_75 B net3 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 net_71 D net_75 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX0 ZN F net_71 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX14 ZN E net_108 VPW NHVT11LL_CKT W=540.00n L=40.00n
XX13 ZN F VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX12 net_108 D VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX10 net_108 C net_100 VPW NHVT11LL_CKT W=540.00n L=40.00n
XX9 net_100 B VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX8 net_100 A1 net4 VPW NHVT11LL_CKT W=540.00n L=40.00n
XX7 net4 A2 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
.ENDS AOAOAOI211111V2_12TH40
.SUBCKT AOAOAOI211111V4_12TH40 A1 A2 B C D E F ZN VDD VSS
XX14 ZN E net_21 VPW NHVT11LL_CKT W=1.08u L=40.00n
XX13 ZN F VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX12 net_21 D VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX10 net_21 C net_29 VPW NHVT11LL_CKT W=1.08u L=40.00n
XX9 net_29 B VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX8 net_29 A1 net4 VPW NHVT11LL_CKT W=1.08u L=40.00n
XX7 net4 A2 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX6 net_64 E VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX5 net_60 C VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX4 net3 A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX3 net3 A1 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX2 net_60 B net3 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 net_64 D net_60 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 ZN F net_64 VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS AOAOAOI211111V4_12TH40
.SUBCKT AOAOAOI211111V8_12TH40 A1 A2 B C D E F ZN VDD VSS
XX14 ZN E net_21 VPW NHVT11LL_CKT W=2.16u L=40.00n
XX13 ZN F VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX12 net_21 D VSS VPW NHVT11LL_CKT W=1.52u L=40.00n
XX10 net_21 C net_29 VPW NHVT11LL_CKT W=2.16u L=40.00n
XX9 net_29 B VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX8 net_29 A1 net4 VPW NHVT11LL_CKT W=2.16u L=40.00n
XX7 net4 A2 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX6 net_64 E VDD VNW PHVT11LL_CKT W=1.72u L=40.00n
XX5 net_60 C VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX4 net3 A2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX3 net3 A1 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX2 net_60 B net3 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 net_64 D net_60 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX0 ZN F net_64 VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS AOAOAOI211111V8_12TH40
.SUBCKT AOAOI2111V1_12TH40 A1 A2 B C D ZN VDD VSS
XX10 net4 A2 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX9 net_11 A1 net4 VPW NHVT11LL_CKT W=380.00n L=40.00n
XX8 net_11 B VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX7 ZN D VSS VPW NHVT11LL_CKT W=190.00n L=40.00n
XX6 ZN C net_11 VPW NHVT11LL_CKT W=380.00n L=40.00n
XX5 ZN D net_30 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX4 net_30 B net3 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX2 net_30 C VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
XX1 net3 A2 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX0 net3 A1 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
.ENDS AOAOI2111V1_12TH40
.SUBCKT AOAOI2111V2_12TH40 A1 A2 B C D ZN VDD VSS
XX10 net4 A2 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX9 net_11 A1 net4 VPW NHVT11LL_CKT W=540.00n L=40.00n
XX8 net_11 B VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX7 ZN D VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX6 ZN C net_11 VPW NHVT11LL_CKT W=540.00n L=40.00n
XX5 ZN D net_30 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX4 net_30 B net3 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX2 net_30 C VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX1 net3 A2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX0 net3 A1 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS AOAOI2111V2_12TH40
.SUBCKT AOAOI2111V4_12TH40 A1 A2 B C D ZN VDD VSS
XX10 net4 A2 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX9 net_11 A1 net4 VPW NHVT11LL_CKT W=1.08u L=40.00n
XX8 net_11 B VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX7 ZN D VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX6 ZN C net_11 VPW NHVT11LL_CKT W=1.08u L=40.00n
XX5 ZN D net_30 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX4 net_30 B net3 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX2 net_30 C VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX1 net3 A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 net3 A1 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS AOAOI2111V4_12TH40
.SUBCKT AOAOI2111V8_12TH40 A1 A2 B C D ZN VDD VSS
XX10 net4 A2 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX9 net_11 A1 net4 VPW NHVT11LL_CKT W=2.16u L=40.00n
XX8 net_11 B VSS VPW NHVT11LL_CKT W=1.52u L=40.00n
XX7 ZN D VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX6 ZN C net_11 VPW NHVT11LL_CKT W=2.16u L=40.00n
XX5 ZN D net_30 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX4 net_30 B net3 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX2 net_30 C VDD VNW PHVT11LL_CKT W=1.72u L=40.00n
XX1 net3 A2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX0 net3 A1 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS AOAOI2111V8_12TH40
.SUBCKT AOI211V0_12TH40 A1 A2 B C ZN VDD VSS
XX4 ZN C VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX3 ZN B VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX9 ZN A1 net18 VPW NHVT11LL_CKT W=0.21u L=40.00n
XX8 net18 A2 VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX2 ZN C net25 VNW PHVT11LL_CKT W=0.365u L=40.00n
XX1 net25 B net34 VNW PHVT11LL_CKT W=0.365u L=40.00n
XX0 net34 A2 VDD VNW PHVT11LL_CKT W=0.365u L=40.00n
XX28 net34 A1 VDD VNW PHVT11LL_CKT W=0.365u L=40.00n
.ENDS AOI211V0_12TH40
.SUBCKT AOI211V1_12TH40 A1 A2 B C ZN VDD VSS
XX4 ZN C VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX3 ZN B VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX9 ZN A1 net18 VPW NHVT11LL_CKT W=0.245u L=40.00n
XX8 net18 A2 VSS VPW NHVT11LL_CKT W=0.245u L=40.00n
XX2 ZN C net25 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX1 net25 B net34 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX0 net34 A2 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX28 net34 A1 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
.ENDS AOI211V1_12TH40
.SUBCKT AOI211V2_12TH40 A1 A2 B C ZN VDD VSS
XX4 ZN C VSS VPW NHVT11LL_CKT W=200.00n L=40.00n
XX3 ZN B VSS VPW NHVT11LL_CKT W=200.00n L=40.00n
XX9 ZN A1 net18 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX8 net18 A2 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX2 ZN C net25 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 net25 B net34 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX0 net34 A2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX28 net34 A1 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS AOI211V2_12TH40
.SUBCKT AOI211V3_12TH40 A1 A2 B C ZN VDD VSS
XX4 ZN C VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX3 ZN B VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX9 ZN A1 net18 VPW NHVT11LL_CKT W=0.49u L=40.00n
XX8 net18 A2 VSS VPW NHVT11LL_CKT W=0.49u L=40.00n
XX2 ZN C net25 VNW PHVT11LL_CKT W=0.86u L=40.00n
XX1 net25 B net34 VNW PHVT11LL_CKT W=0.86u L=40.00n
XX0 net34 A2 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX28 net34 A1 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
.ENDS AOI211V3_12TH40
.SUBCKT AOI211V4_12TH40 A1 A2 B C ZN VDD VSS
XX4 ZN C VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX3 ZN B VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX9 ZN A1 net18 VPW NHVT11LL_CKT W=0.7u L=40.00n
XX8 net18 A2 VSS VPW NHVT11LL_CKT W=0.7u L=40.00n
XX2 ZN C net25 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 net25 B net34 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 net34 A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX28 net34 A1 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS AOI211V4_12TH40
.SUBCKT AOI211V6_12TH40 A1 A2 B C ZN VDD VSS
XX4 ZN C VSS VPW NHVT11LL_CKT W=0.6u L=40.00n
XX3 ZN B VSS VPW NHVT11LL_CKT W=0.6u L=40.00n
XX9 ZN A1 net18 VPW NHVT11LL_CKT W=1.05u L=40.00n
XX8 net18 A2 VSS VPW NHVT11LL_CKT W=1.05u L=40.00n
XX2 ZN C net25 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX1 net25 B net34 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX0 net34 A2 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX28 net34 A1 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS AOI211V6_12TH40
.SUBCKT AOI211V8_12TH40 A1 A2 B C ZN VDD VSS
XX4 ZN C VSS VPW NHVT11LL_CKT W=0.8u L=40.00n
XX3 ZN B VSS VPW NHVT11LL_CKT W=0.8u L=40.00n
XX9 ZN A1 net18 VPW NHVT11LL_CKT W=1.4u L=40.00n
XX8 net18 A2 VSS VPW NHVT11LL_CKT W=1.4u L=40.00n
XX2 ZN C net25 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 net25 B net34 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX0 net34 A2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX28 net34 A1 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS AOI211V8_12TH40
.SUBCKT AOI21BV0_12TH40 A B1 B2 ZN VDD VSS
XX3 net21 A VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX2 ZN net21 VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX9 ZN B1 net33 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX8 net33 B2 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX4 net21 A VDD VNW PHVT11LL_CKT W=0.135u L=40.00n
XX1 ZN net21 net17 VNW PHVT11LL_CKT W=0.305u L=40.00n
XX0 net17 B2 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX28 net17 B1 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
.ENDS AOI21BV0_12TH40
.SUBCKT AOI21BV12_12TH40 A B1 B2 ZN VDD VSS
XX3 net21 A VSS VPW NHVT11LL_CKT W=0.72u L=40.00n
XX2 ZN net21 VSS VPW NHVT11LL_CKT W=1.71u L=40.00n
XX9 ZN B1 net33 VPW NHVT11LL_CKT W=3.03u L=40.00n
XX8 net33 B2 VSS VPW NHVT11LL_CKT W=3.03u L=40.00n
XX4 net21 A VDD VNW PHVT11LL_CKT W=0.82u L=40.00n
XX1 ZN net21 net17 VNW PHVT11LL_CKT W=3.66u L=40.00n
XX0 net17 B2 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX28 net17 B1 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
.ENDS AOI21BV12_12TH40
.SUBCKT AOI21BV16_12TH40 A B1 B2 ZN VDD VSS
XX3 net21 A VSS VPW NHVT11LL_CKT W=0.95u L=40.00n
XX2 ZN net21 VSS VPW NHVT11LL_CKT W=2.28u L=40.00n
XX9 ZN B1 net33 VPW NHVT11LL_CKT W=4.04u L=40.00n
XX8 net33 B2 VSS VPW NHVT11LL_CKT W=4.04u L=40.00n
XX4 net21 A VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX1 ZN net21 net17 VNW PHVT11LL_CKT W=4.88u L=40.00n
XX0 net17 B2 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX28 net17 B1 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
.ENDS AOI21BV16_12TH40
.SUBCKT AOI21BV1_12TH40 A B1 B2 ZN VDD VSS
XX3 net21 A VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX2 ZN net21 VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX9 ZN B1 net33 VPW NHVT11LL_CKT W=0.355u L=40.00n
XX8 net33 B2 VSS VPW NHVT11LL_CKT W=0.355u L=40.00n
XX4 net21 A VDD VNW PHVT11LL_CKT W=0.135u L=40.00n
XX1 ZN net21 net17 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX0 net17 B2 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX28 net17 B1 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
.ENDS AOI21BV1_12TH40
.SUBCKT AOI21BV2_12TH40 A B1 B2 ZN VDD VSS
XX3 net21 A VSS VPW NHVT11LL_CKT W=145.00n L=40.00n
XX2 ZN net21 VSS VPW NHVT11LL_CKT W=285.00n L=40.00n
XX9 ZN B1 net33 VPW NHVT11LL_CKT W=505.00n L=40.00n
XX8 net33 B2 VSS VPW NHVT11LL_CKT W=505.00n L=40.00n
XX4 net21 A VDD VNW PHVT11LL_CKT W=165.00n L=40.00n
XX1 ZN net21 net17 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX0 net17 B2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX28 net17 B1 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS AOI21BV2_12TH40
.SUBCKT AOI21BV3_12TH40 A B1 B2 ZN VDD VSS
XX3 net21 A VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX2 ZN net21 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX9 ZN B1 net33 VPW NHVT11LL_CKT W=0.71u L=40.00n
XX8 net33 B2 VSS VPW NHVT11LL_CKT W=0.71u L=40.00n
XX4 net21 A VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX1 ZN net21 net17 VNW PHVT11LL_CKT W=0.86u L=40.00n
XX0 net17 B2 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX28 net17 B1 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
.ENDS AOI21BV3_12TH40
.SUBCKT AOI21BV4_12TH40 A B1 B2 ZN VDD VSS
XX3 net21 A VSS VPW NHVT11LL_CKT W=0.255u L=40.00n
XX2 ZN net21 VSS VPW NHVT11LL_CKT W=0.57u L=40.00n
XX9 ZN B1 net33 VPW NHVT11LL_CKT W=1.01u L=40.00n
XX8 net33 B2 VSS VPW NHVT11LL_CKT W=1.01u L=40.00n
XX4 net21 A VDD VNW PHVT11LL_CKT W=0.29u L=40.00n
XX1 ZN net21 net17 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 net17 B2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX28 net17 B1 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS AOI21BV4_12TH40
.SUBCKT AOI21BV6_12TH40 A B1 B2 ZN VDD VSS
XX3 net21 A VSS VPW NHVT11LL_CKT W=0.365u L=40.00n
XX2 ZN net21 VSS VPW NHVT11LL_CKT W=0.855u L=40.00n
XX9 ZN B1 net33 VPW NHVT11LL_CKT W=1.515u L=40.00n
XX8 net33 B2 VSS VPW NHVT11LL_CKT W=1.515u L=40.00n
XX4 net21 A VDD VNW PHVT11LL_CKT W=0.415u L=40.00n
XX1 ZN net21 net17 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX0 net17 B2 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX28 net17 B1 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS AOI21BV6_12TH40
.SUBCKT AOI21BV8_12TH40 A B1 B2 ZN VDD VSS
XX3 net21 A VSS VPW NHVT11LL_CKT W=0.48u L=40.00n
XX2 ZN net21 VSS VPW NHVT11LL_CKT W=1.14u L=40.00n
XX9 ZN B1 net33 VPW NHVT11LL_CKT W=2.02u L=40.00n
XX8 net33 B2 VSS VPW NHVT11LL_CKT W=2.02u L=40.00n
XX4 net21 A VDD VNW PHVT11LL_CKT W=0.545u L=40.00n
XX1 ZN net21 net17 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX0 net17 B2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX28 net17 B1 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS AOI21BV8_12TH40
.SUBCKT AOI21V0_12TH40 A1 A2 B ZN VDD VSS
XX8 net5 A2 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX9 ZN A1 net5 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX2 ZN B VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX28 net17 A1 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX0 net17 A2 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX1 ZN B net17 VNW PHVT11LL_CKT W=0.305u L=40.00n
.ENDS AOI21V0_12TH40
.SUBCKT AOI21V12_12TH40 A1 A2 B ZN VDD VSS
XX8 net5 A2 VSS VPW NHVT11LL_CKT W=3.03u L=40.00n
XX9 ZN A1 net5 VPW NHVT11LL_CKT W=3.03u L=40.00n
XX2 ZN B VSS VPW NHVT11LL_CKT W=1.71u L=40.00n
XX28 net17 A1 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX0 net17 A2 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX1 ZN B net17 VNW PHVT11LL_CKT W=3.66u L=40.00n
.ENDS AOI21V12_12TH40
.SUBCKT AOI21V16_12TH40 A1 A2 B ZN VDD VSS
XX8 net5 A2 VSS VPW NHVT11LL_CKT W=4.04u L=40.00n
XX9 ZN A1 net5 VPW NHVT11LL_CKT W=4.04u L=40.00n
XX2 ZN B VSS VPW NHVT11LL_CKT W=2.28u L=40.00n
XX28 net17 A1 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX0 net17 A2 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX1 ZN B net17 VNW PHVT11LL_CKT W=4.88u L=40.00n
.ENDS AOI21V16_12TH40
.SUBCKT AOI21V1_12TH40 A1 A2 B ZN VDD VSS
XX8 net5 A2 VSS VPW NHVT11LL_CKT W=0.355u L=40.00n
XX9 ZN A1 net5 VPW NHVT11LL_CKT W=0.355u L=40.00n
XX2 ZN B VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX28 net17 A1 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX0 net17 A2 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX1 ZN B net17 VNW PHVT11LL_CKT W=0.43u L=40.00n
.ENDS AOI21V1_12TH40
.SUBCKT AOI21V2_12TH40 A1 A2 B ZN VDD VSS
XX8 net5 A2 VSS VPW NHVT11LL_CKT W=505.00n L=40.00n
XX9 ZN A1 net5 VPW NHVT11LL_CKT W=505.00n L=40.00n
XX2 ZN B VSS VPW NHVT11LL_CKT W=285.00n L=40.00n
XX28 net17 A1 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX0 net17 A2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 ZN B net17 VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS AOI21V2_12TH40
.SUBCKT AOI21V3_12TH40 A1 A2 B ZN VDD VSS
XX8 net5 A2 VSS VPW NHVT11LL_CKT W=0.71u L=40.00n
XX9 ZN A1 net5 VPW NHVT11LL_CKT W=0.71u L=40.00n
XX2 ZN B VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX28 net17 A1 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX0 net17 A2 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX1 ZN B net17 VNW PHVT11LL_CKT W=0.86u L=40.00n
.ENDS AOI21V3_12TH40
.SUBCKT AOI21V4_12TH40 A1 A2 B ZN VDD VSS
XX8 net5 A2 VSS VPW NHVT11LL_CKT W=1.01u L=40.00n
XX9 ZN A1 net5 VPW NHVT11LL_CKT W=1.01u L=40.00n
XX2 ZN B VSS VPW NHVT11LL_CKT W=0.57u L=40.00n
XX28 net17 A1 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 net17 A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 ZN B net17 VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS AOI21V4_12TH40
.SUBCKT AOI21V6_12TH40 A1 A2 B ZN VDD VSS
XX8 net5 A2 VSS VPW NHVT11LL_CKT W=1.515u L=40.00n
XX9 ZN A1 net5 VPW NHVT11LL_CKT W=1.515u L=40.00n
XX2 ZN B VSS VPW NHVT11LL_CKT W=0.855u L=40.00n
XX28 net17 A1 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX0 net17 A2 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX1 ZN B net17 VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS AOI21V6_12TH40
.SUBCKT AOI21V8_12TH40 A1 A2 B ZN VDD VSS
XX8 net5 A2 VSS VPW NHVT11LL_CKT W=2.02u L=40.00n
XX9 ZN A1 net5 VPW NHVT11LL_CKT W=2.02u L=40.00n
XX2 ZN B VSS VPW NHVT11LL_CKT W=1.14u L=40.00n
XX28 net17 A1 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX0 net17 A2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 ZN B net17 VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS AOI21V8_12TH40
.SUBCKT AOI221V0_12TH40 A1 A2 B1 B2 C ZN VDD VSS
XX4 ZN C VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX2 ZN B1 net31 VPW NHVT11LL_CKT W=0.21u L=40.00n
XX9 ZN A1 net43 VPW NHVT11LL_CKT W=0.21u L=40.00n
XX8 net43 A2 VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX3 net31 B2 VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX6 net26 A1 VDD VNW PHVT11LL_CKT W=0.365u L=40.00n
XX5 net26 A2 VDD VNW PHVT11LL_CKT W=0.365u L=40.00n
XX1 ZN C net23 VNW PHVT11LL_CKT W=0.365u L=40.00n
XX0 net23 B2 net26 VNW PHVT11LL_CKT W=0.365u L=40.00n
XX28 net23 B1 net26 VNW PHVT11LL_CKT W=0.365u L=40.00n
.ENDS AOI221V0_12TH40
.SUBCKT AOI221V1_12TH40 A1 A2 B1 B2 C ZN VDD VSS
XX4 ZN C VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX2 ZN B1 net31 VPW NHVT11LL_CKT W=0.245u L=40.00n
XX9 ZN A1 net43 VPW NHVT11LL_CKT W=0.245u L=40.00n
XX8 net43 A2 VSS VPW NHVT11LL_CKT W=0.245u L=40.00n
XX3 net31 B2 VSS VPW NHVT11LL_CKT W=0.245u L=40.00n
XX6 net26 A1 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX5 net26 A2 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX1 ZN C net23 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX0 net23 B2 net26 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX28 net23 B1 net26 VNW PHVT11LL_CKT W=0.43u L=40.00n
.ENDS AOI221V1_12TH40
.SUBCKT AOI221V2_12TH40 A1 A2 B1 B2 C ZN VDD VSS
XX4 ZN C VSS VPW NHVT11LL_CKT W=200.00n L=40.00n
XX2 ZN B1 net31 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX9 ZN A1 net43 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX8 net43 A2 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX3 net31 B2 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX6 net26 A1 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX5 net26 A2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 ZN C net23 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX0 net23 B2 net26 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX28 net23 B1 net26 VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS AOI221V2_12TH40
.SUBCKT AOI221V3_12TH40 A1 A2 B1 B2 C ZN VDD VSS
XX4 ZN C VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX2 ZN B1 net31 VPW NHVT11LL_CKT W=0.49u L=40.00n
XX9 ZN A1 net43 VPW NHVT11LL_CKT W=0.49u L=40.00n
XX8 net43 A2 VSS VPW NHVT11LL_CKT W=0.49u L=40.00n
XX3 net31 B2 VSS VPW NHVT11LL_CKT W=0.49u L=40.00n
XX6 net26 A1 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX5 net26 A2 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX1 ZN C net23 VNW PHVT11LL_CKT W=0.86u L=40.00n
XX0 net23 B2 net26 VNW PHVT11LL_CKT W=0.86u L=40.00n
XX28 net23 B1 net26 VNW PHVT11LL_CKT W=0.86u L=40.00n
.ENDS AOI221V3_12TH40
.SUBCKT AOI221V4_12TH40 A1 A2 B1 B2 C ZN VDD VSS
XX4 ZN C VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX2 ZN B1 net31 VPW NHVT11LL_CKT W=0.7u L=40.00n
XX9 ZN A1 net43 VPW NHVT11LL_CKT W=0.7u L=40.00n
XX8 net43 A2 VSS VPW NHVT11LL_CKT W=0.7u L=40.00n
XX3 net31 B2 VSS VPW NHVT11LL_CKT W=0.7u L=40.00n
XX6 net26 A1 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX5 net26 A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 ZN C net23 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 net23 B2 net26 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX28 net23 B1 net26 VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS AOI221V4_12TH40
.SUBCKT AOI221V6_12TH40 A1 A2 B1 B2 C ZN VDD VSS
XX4 ZN C VSS VPW NHVT11LL_CKT W=0.6u L=40.00n
XX2 ZN B1 net31 VPW NHVT11LL_CKT W=1.05u L=40.00n
XX9 ZN A1 net43 VPW NHVT11LL_CKT W=1.05u L=40.00n
XX8 net43 A2 VSS VPW NHVT11LL_CKT W=1.05u L=40.00n
XX3 net31 B2 VSS VPW NHVT11LL_CKT W=1.05u L=40.00n
XX6 net26 A1 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX5 net26 A2 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX1 ZN C net23 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX0 net23 B2 net26 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX28 net23 B1 net26 VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS AOI221V6_12TH40
.SUBCKT AOI221V8_12TH40 A1 A2 B1 B2 C ZN VDD VSS
XX4 ZN C VSS VPW NHVT11LL_CKT W=0.8u L=40.00n
XX2 ZN B1 net31 VPW NHVT11LL_CKT W=1.4u L=40.00n
XX9 ZN A1 net43 VPW NHVT11LL_CKT W=1.4u L=40.00n
XX8 net43 A2 VSS VPW NHVT11LL_CKT W=1.4u L=40.00n
XX3 net31 B2 VSS VPW NHVT11LL_CKT W=1.4u L=40.00n
XX6 net26 A1 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX5 net26 A2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 ZN C net23 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX0 net23 B2 net26 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX28 net23 B1 net26 VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS AOI221V8_12TH40
.SUBCKT AOI222V0_12TH40 A1 A2 B1 B2 C1 C2 ZN VDD VSS
XX7 net8 C2 VSS VPW NHVT11LL_CKT W=0.175u L=40.00n
XX3 net12 B2 VSS VPW NHVT11LL_CKT W=0.175u L=40.00n
XX8 net16 A2 VSS VPW NHVT11LL_CKT W=0.175u L=40.00n
XX9 ZN A1 net16 VPW NHVT11LL_CKT W=0.175u L=40.00n
XX2 ZN B1 net12 VPW NHVT11LL_CKT W=0.175u L=40.00n
XX4 ZN C1 net8 VPW NHVT11LL_CKT W=0.175u L=40.00n
XX10 ZN C2 net39 VNW PHVT11LL_CKT W=0.305u L=40.00n
XX28 net39 B1 net43 VNW PHVT11LL_CKT W=0.305u L=40.00n
XX0 net39 B2 net43 VNW PHVT11LL_CKT W=0.305u L=40.00n
XX1 ZN C1 net39 VNW PHVT11LL_CKT W=0.305u L=40.00n
XX5 net43 A2 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX6 net43 A1 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
.ENDS AOI222V0_12TH40
.SUBCKT AOI222V1_12TH40 A1 A2 B1 B2 C1 C2 ZN VDD VSS
XX7 net8 C2 VSS VPW NHVT11LL_CKT W=0.245u L=40.00n
XX3 net12 B2 VSS VPW NHVT11LL_CKT W=0.245u L=40.00n
XX8 net16 A2 VSS VPW NHVT11LL_CKT W=0.245u L=40.00n
XX9 ZN A1 net16 VPW NHVT11LL_CKT W=0.245u L=40.00n
XX2 ZN B1 net12 VPW NHVT11LL_CKT W=0.245u L=40.00n
XX4 ZN C1 net8 VPW NHVT11LL_CKT W=0.245u L=40.00n
XX10 ZN C2 net39 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX28 net39 B1 net43 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX0 net39 B2 net43 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX1 ZN C1 net39 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX5 net43 A2 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX6 net43 A1 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
.ENDS AOI222V1_12TH40
.SUBCKT AOI222V2_12TH40 A1 A2 B1 B2 C1 C2 ZN VDD VSS
XX7 net8 C2 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX3 net12 B2 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX8 net16 A2 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX9 ZN A1 net16 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX2 ZN B1 net12 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX4 ZN C1 net8 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX10 ZN C2 net39 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX28 net39 B1 net43 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX0 net39 B2 net43 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 ZN C1 net39 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX5 net43 A2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX6 net43 A1 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS AOI222V2_12TH40
.SUBCKT AOI222V3_12TH40 A1 A2 B1 B2 C1 C2 ZN VDD VSS
XX7 net8 C2 VSS VPW NHVT11LL_CKT W=0.49u L=40.00n
XX3 net12 B2 VSS VPW NHVT11LL_CKT W=0.49u L=40.00n
XX8 net16 A2 VSS VPW NHVT11LL_CKT W=0.49u L=40.00n
XX9 ZN A1 net16 VPW NHVT11LL_CKT W=0.49u L=40.00n
XX2 ZN B1 net12 VPW NHVT11LL_CKT W=0.49u L=40.00n
XX4 ZN C1 net8 VPW NHVT11LL_CKT W=0.49u L=40.00n
XX10 ZN C2 net39 VNW PHVT11LL_CKT W=0.86u L=40.00n
XX28 net39 B1 net43 VNW PHVT11LL_CKT W=0.86u L=40.00n
XX0 net39 B2 net43 VNW PHVT11LL_CKT W=0.86u L=40.00n
XX1 ZN C1 net39 VNW PHVT11LL_CKT W=0.86u L=40.00n
XX5 net43 A2 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX6 net43 A1 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
.ENDS AOI222V3_12TH40
.SUBCKT AOI222V4_12TH40 A1 A2 B1 B2 C1 C2 ZN VDD VSS
XX7 net8 C2 VSS VPW NHVT11LL_CKT W=0.7u L=40.00n
XX3 net12 B2 VSS VPW NHVT11LL_CKT W=0.7u L=40.00n
XX8 net16 A2 VSS VPW NHVT11LL_CKT W=0.7u L=40.00n
XX9 ZN A1 net16 VPW NHVT11LL_CKT W=0.7u L=40.00n
XX2 ZN B1 net12 VPW NHVT11LL_CKT W=0.7u L=40.00n
XX4 ZN C1 net8 VPW NHVT11LL_CKT W=0.7u L=40.00n
XX10 ZN C2 net39 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX28 net39 B1 net43 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 net39 B2 net43 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 ZN C1 net39 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX5 net43 A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX6 net43 A1 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS AOI222V4_12TH40
.SUBCKT AOI222V6_12TH40 A1 A2 B1 B2 C1 C2 ZN VDD VSS
XX7 net8 C2 VSS VPW NHVT11LL_CKT W=1.05u L=40.00n
XX3 net12 B2 VSS VPW NHVT11LL_CKT W=1.05u L=40.00n
XX8 net16 A2 VSS VPW NHVT11LL_CKT W=1.05u L=40.00n
XX9 ZN A1 net16 VPW NHVT11LL_CKT W=1.05u L=40.00n
XX2 ZN B1 net12 VPW NHVT11LL_CKT W=1.05u L=40.00n
XX4 ZN C1 net8 VPW NHVT11LL_CKT W=1.05u L=40.00n
XX10 ZN C2 net39 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX28 net39 B1 net43 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX0 net39 B2 net43 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX1 ZN C1 net39 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX5 net43 A2 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX6 net43 A1 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS AOI222V6_12TH40
.SUBCKT AOI222V8_12TH40 A1 A2 B1 B2 C1 C2 ZN VDD VSS
XX7 net8 C2 VSS VPW NHVT11LL_CKT W=1.4u L=40.00n
XX3 net12 B2 VSS VPW NHVT11LL_CKT W=1.4u L=40.00n
XX8 net16 A2 VSS VPW NHVT11LL_CKT W=1.4u L=40.00n
XX9 ZN A1 net16 VPW NHVT11LL_CKT W=1.4u L=40.00n
XX2 ZN B1 net12 VPW NHVT11LL_CKT W=1.4u L=40.00n
XX4 ZN C1 net8 VPW NHVT11LL_CKT W=1.4u L=40.00n
XX10 ZN C2 net39 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX28 net39 B1 net43 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX0 net39 B2 net43 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 ZN C1 net39 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX5 net43 A2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX6 net43 A1 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS AOI222V8_12TH40
.SUBCKT AOI22BBV0_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX20 net34 B2 VSS VPW NHVT11LL_CKT W=0.205u L=40.00n
XX19 ZN B1 net34 VPW NHVT11LL_CKT W=0.205u L=40.00n
XX18 ZN net30 VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX14 net30 A1 VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX13 net30 A2 VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX17 ZN net30 net22 VNW PHVT11LL_CKT W=0.305u L=40.00n
XX16 net22 B2 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX15 net22 B1 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX12 net30 A1 net9 VNW PHVT11LL_CKT W=0.215u L=40.00n
XX11 net9 A2 VDD VNW PHVT11LL_CKT W=0.215u L=40.00n
.ENDS AOI22BBV0_12TH40
.SUBCKT AOI22BBV12_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX20 net34 B2 VSS VPW NHVT11LL_CKT W=3.03u L=40.00n
XX19 ZN B1 net34 VPW NHVT11LL_CKT W=3.03u L=40.00n
XX18 ZN net30 VSS VPW NHVT11LL_CKT W=1.71u L=40.00n
XX14 net30 A1 VSS VPW NHVT11LL_CKT W=1.095u L=40.00n
XX13 net30 A2 VSS VPW NHVT11LL_CKT W=1.095u L=40.00n
XX17 ZN net30 net22 VNW PHVT11LL_CKT W=3.66u L=40.00n
XX16 net22 B2 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX15 net22 B1 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX12 net30 A1 net9 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX11 net9 A2 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS AOI22BBV12_12TH40
.SUBCKT AOI22BBV16_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX20 net34 B2 VSS VPW NHVT11LL_CKT W=4.04u L=40.00n
XX19 ZN B1 net34 VPW NHVT11LL_CKT W=4.04u L=40.00n
XX18 ZN net30 VSS VPW NHVT11LL_CKT W=2.28u L=40.00n
XX14 net30 A1 VSS VPW NHVT11LL_CKT W=1.46u L=40.00n
XX13 net30 A2 VSS VPW NHVT11LL_CKT W=1.46u L=40.00n
XX17 ZN net30 net22 VNW PHVT11LL_CKT W=4.88u L=40.00n
XX16 net22 B2 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX15 net22 B1 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX12 net30 A1 net9 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX11 net9 A2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS AOI22BBV16_12TH40
.SUBCKT AOI22BBV1_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX20 net34 B2 VSS VPW NHVT11LL_CKT W=0.355u L=40.00n
XX19 ZN B1 net34 VPW NHVT11LL_CKT W=0.355u L=40.00n
XX18 ZN net30 VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX14 net30 A1 VSS VPW NHVT11LL_CKT W=0.165u L=40.00n
XX13 net30 A2 VSS VPW NHVT11LL_CKT W=0.165u L=40.00n
XX17 ZN net30 net22 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX16 net22 B2 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX15 net22 B1 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX12 net30 A1 net9 VNW PHVT11LL_CKT W=0.28u L=40.00n
XX11 net9 A2 VDD VNW PHVT11LL_CKT W=0.28u L=40.00n
.ENDS AOI22BBV1_12TH40
.SUBCKT AOI22BBV2_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX20 net34 B2 VSS VPW NHVT11LL_CKT W=505.00n L=40.00n
XX19 ZN B1 net34 VPW NHVT11LL_CKT W=505.00n L=40.00n
XX18 ZN net30 VSS VPW NHVT11LL_CKT W=285.00n L=40.00n
XX14 net30 A1 VSS VPW NHVT11LL_CKT W=210.00n L=40.00n
XX13 net30 A2 VSS VPW NHVT11LL_CKT W=210.00n L=40.00n
XX17 ZN net30 net22 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX16 net22 B2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX15 net22 B1 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX12 net30 A1 net9 VNW PHVT11LL_CKT W=345.00n L=40.00n
XX11 net9 A2 VDD VNW PHVT11LL_CKT W=345.00n L=40.00n
.ENDS AOI22BBV2_12TH40
.SUBCKT AOI22BBV3_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX20 net34 B2 VSS VPW NHVT11LL_CKT W=0.71u L=40.00n
XX19 ZN B1 net34 VPW NHVT11LL_CKT W=0.71u L=40.00n
XX18 ZN net30 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX14 net30 A1 VSS VPW NHVT11LL_CKT W=0.275u L=40.00n
XX13 net30 A2 VSS VPW NHVT11LL_CKT W=0.275u L=40.00n
XX17 ZN net30 net22 VNW PHVT11LL_CKT W=0.86u L=40.00n
XX16 net22 B2 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX15 net22 B1 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX12 net30 A1 net9 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX11 net9 A2 VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
.ENDS AOI22BBV3_12TH40
.SUBCKT AOI22BBV4_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX20 net34 B2 VSS VPW NHVT11LL_CKT W=1.01u L=40.00n
XX19 ZN B1 net34 VPW NHVT11LL_CKT W=1.01u L=40.00n
XX18 ZN net30 VSS VPW NHVT11LL_CKT W=0.57u L=40.00n
XX14 net30 A1 VSS VPW NHVT11LL_CKT W=0.365u L=40.00n
XX13 net30 A2 VSS VPW NHVT11LL_CKT W=0.365u L=40.00n
XX17 ZN net30 net22 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX16 net22 B2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX15 net22 B1 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX12 net30 A1 net9 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX11 net9 A2 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
.ENDS AOI22BBV4_12TH40
.SUBCKT AOI22BBV6_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX20 net34 B2 VSS VPW NHVT11LL_CKT W=1.515u L=40.00n
XX19 ZN B1 net34 VPW NHVT11LL_CKT W=1.515u L=40.00n
XX18 ZN net30 VSS VPW NHVT11LL_CKT W=0.855u L=40.00n
XX14 net30 A1 VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX13 net30 A2 VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX17 ZN net30 net22 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX16 net22 B2 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX15 net22 B1 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX12 net30 A1 net9 VNW PHVT11LL_CKT W=0.9u L=40.00n
XX11 net9 A2 VDD VNW PHVT11LL_CKT W=0.9u L=40.00n
.ENDS AOI22BBV6_12TH40
.SUBCKT AOI22BBV8_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX20 net34 B2 VSS VPW NHVT11LL_CKT W=2.02u L=40.00n
XX19 ZN B1 net34 VPW NHVT11LL_CKT W=2.02u L=40.00n
XX18 ZN net30 VSS VPW NHVT11LL_CKT W=1.14u L=40.00n
XX14 net30 A1 VSS VPW NHVT11LL_CKT W=0.73u L=40.00n
XX13 net30 A2 VSS VPW NHVT11LL_CKT W=0.73u L=40.00n
XX17 ZN net30 net22 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX16 net22 B2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX15 net22 B1 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX12 net30 A1 net9 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX11 net9 A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS AOI22BBV8_12TH40
.SUBCKT AOI22V0_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX8 net22 A2 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX9 ZN A1 net22 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX3 ZN B1 net34 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX4 net34 B2 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX28 net17 A1 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX0 net17 A2 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX1 ZN B1 net17 VNW PHVT11LL_CKT W=0.305u L=40.00n
XX2 ZN B2 net17 VNW PHVT11LL_CKT W=0.305u L=40.00n
.ENDS AOI22V0_12TH40
.SUBCKT AOI22V12_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX8 net22 A2 VSS VPW NHVT11LL_CKT W=3.03u L=40.00n
XX9 ZN A1 net22 VPW NHVT11LL_CKT W=3.03u L=40.00n
XX3 ZN B1 net34 VPW NHVT11LL_CKT W=3.03u L=40.00n
XX4 net34 B2 VSS VPW NHVT11LL_CKT W=3.03u L=40.00n
XX28 net17 A1 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX0 net17 A2 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX1 ZN B1 net17 VNW PHVT11LL_CKT W=3.66u L=40.00n
XX2 ZN B2 net17 VNW PHVT11LL_CKT W=3.66u L=40.00n
.ENDS AOI22V12_12TH40
.SUBCKT AOI22V16_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX8 net22 A2 VSS VPW NHVT11LL_CKT W=4.04u L=40.00n
XX9 ZN A1 net22 VPW NHVT11LL_CKT W=4.04u L=40.00n
XX3 ZN B1 net34 VPW NHVT11LL_CKT W=4.04u L=40.00n
XX4 net34 B2 VSS VPW NHVT11LL_CKT W=4.04u L=40.00n
XX28 net17 A1 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX0 net17 A2 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX1 ZN B1 net17 VNW PHVT11LL_CKT W=4.88u L=40.00n
XX2 ZN B2 net17 VNW PHVT11LL_CKT W=4.88u L=40.00n
.ENDS AOI22V16_12TH40
.SUBCKT AOI22V1_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX8 net22 A2 VSS VPW NHVT11LL_CKT W=0.355u L=40.00n
XX9 ZN A1 net22 VPW NHVT11LL_CKT W=0.355u L=40.00n
XX3 ZN B1 net34 VPW NHVT11LL_CKT W=0.355u L=40.00n
XX4 net34 B2 VSS VPW NHVT11LL_CKT W=0.355u L=40.00n
XX28 net17 A1 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX0 net17 A2 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX1 ZN B1 net17 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX2 ZN B2 net17 VNW PHVT11LL_CKT W=0.43u L=40.00n
.ENDS AOI22V1_12TH40
.SUBCKT AOI22V2_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX8 net22 A2 VSS VPW NHVT11LL_CKT W=505.00n L=40.00n
XX9 ZN A1 net22 VPW NHVT11LL_CKT W=505.00n L=40.00n
XX3 ZN B1 net34 VPW NHVT11LL_CKT W=505.00n L=40.00n
XX4 net34 B2 VSS VPW NHVT11LL_CKT W=505.00n L=40.00n
XX28 net17 A1 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX0 net17 A2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 ZN B1 net17 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX2 ZN B2 net17 VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS AOI22V2_12TH40
.SUBCKT AOI22V3_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX8 net22 A2 VSS VPW NHVT11LL_CKT W=0.71u L=40.00n
XX9 ZN A1 net22 VPW NHVT11LL_CKT W=0.71u L=40.00n
XX3 ZN B1 net34 VPW NHVT11LL_CKT W=0.71u L=40.00n
XX4 net34 B2 VSS VPW NHVT11LL_CKT W=0.71u L=40.00n
XX28 net17 A1 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX0 net17 A2 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX1 ZN B1 net17 VNW PHVT11LL_CKT W=0.86u L=40.00n
XX2 ZN B2 net17 VNW PHVT11LL_CKT W=0.86u L=40.00n
.ENDS AOI22V3_12TH40
.SUBCKT AOI22V4_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX8 net22 A2 VSS VPW NHVT11LL_CKT W=1.01u L=40.00n
XX9 ZN A1 net22 VPW NHVT11LL_CKT W=1.01u L=40.00n
XX3 ZN B1 net34 VPW NHVT11LL_CKT W=1.01u L=40.00n
XX4 net34 B2 VSS VPW NHVT11LL_CKT W=1.01u L=40.00n
XX28 net17 A1 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 net17 A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 ZN B1 net17 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX2 ZN B2 net17 VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS AOI22V4_12TH40
.SUBCKT AOI22V6_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX8 net22 A2 VSS VPW NHVT11LL_CKT W=1.515u L=40.00n
XX9 ZN A1 net22 VPW NHVT11LL_CKT W=1.515u L=40.00n
XX3 ZN B1 net34 VPW NHVT11LL_CKT W=1.515u L=40.00n
XX4 net34 B2 VSS VPW NHVT11LL_CKT W=1.515u L=40.00n
XX28 net17 A1 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX0 net17 A2 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX1 ZN B1 net17 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX2 ZN B2 net17 VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS AOI22V6_12TH40
.SUBCKT AOI22V8_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX8 net22 A2 VSS VPW NHVT11LL_CKT W=2.02u L=40.00n
XX9 ZN A1 net22 VPW NHVT11LL_CKT W=2.02u L=40.00n
XX3 ZN B1 net34 VPW NHVT11LL_CKT W=2.02u L=40.00n
XX4 net34 B2 VSS VPW NHVT11LL_CKT W=2.02u L=40.00n
XX28 net17 A1 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX0 net17 A2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 ZN B1 net17 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX2 ZN B2 net17 VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS AOI22V8_12TH40
.SUBCKT AOI2XB1V0_12TH40 A B1 B2 ZN VDD VSS
XX4 net21 B2 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX2 ZN A VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX9 ZN B1 net25 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX8 net25 net21 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX3 net21 B2 VDD VNW PHVT11LL_CKT W=0.135u L=40.00n
XX1 ZN A net9 VNW PHVT11LL_CKT W=0.305u L=40.00n
XX0 net9 B1 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX28 net9 net21 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
.ENDS AOI2XB1V0_12TH40
.SUBCKT AOI2XB1V12_12TH40 A B1 B2 ZN VDD VSS
XX4 net21 B2 VSS VPW NHVT11LL_CKT W=0.87u L=40.00n
XX2 ZN A VSS VPW NHVT11LL_CKT W=1.71u L=40.00n
XX9 ZN B1 net25 VPW NHVT11LL_CKT W=3.03u L=40.00n
XX8 net25 net21 VSS VPW NHVT11LL_CKT W=3.03u L=40.00n
XX3 net21 B2 VDD VNW PHVT11LL_CKT W=1u L=40.00n
XX1 ZN A net9 VNW PHVT11LL_CKT W=3.66u L=40.00n
XX0 net9 B1 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX28 net9 net21 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
.ENDS AOI2XB1V12_12TH40
.SUBCKT AOI2XB1V16_12TH40 A B1 B2 ZN VDD VSS
XX4 net21 B2 VSS VPW NHVT11LL_CKT W=1.185u L=40.00n
XX2 ZN A VSS VPW NHVT11LL_CKT W=2.28u L=40.00n
XX9 ZN B1 net25 VPW NHVT11LL_CKT W=4.04u L=40.00n
XX8 net25 net21 VSS VPW NHVT11LL_CKT W=4.04u L=40.00n
XX3 net21 B2 VDD VNW PHVT11LL_CKT W=1.35u L=40.00n
XX1 ZN A net9 VNW PHVT11LL_CKT W=4.88u L=40.00n
XX0 net9 B1 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX28 net9 net21 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
.ENDS AOI2XB1V16_12TH40
.SUBCKT AOI2XB1V1_12TH40 A B1 B2 ZN VDD VSS
XX4 net21 B2 VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX2 ZN A VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX9 ZN B1 net25 VPW NHVT11LL_CKT W=0.355u L=40.00n
XX8 net25 net21 VSS VPW NHVT11LL_CKT W=0.355u L=40.00n
XX3 net21 B2 VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX1 ZN A net9 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX0 net9 B1 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX28 net9 net21 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
.ENDS AOI2XB1V1_12TH40
.SUBCKT AOI2XB1V2_12TH40 A B1 B2 ZN VDD VSS
XX4 net21 B2 VSS VPW NHVT11LL_CKT W=170.00n L=40.00n
XX2 ZN A VSS VPW NHVT11LL_CKT W=285.00n L=40.00n
XX9 ZN B1 net25 VPW NHVT11LL_CKT W=505.00n L=40.00n
XX8 net25 net21 VSS VPW NHVT11LL_CKT W=505.00n L=40.00n
XX3 net21 B2 VDD VNW PHVT11LL_CKT W=195.00n L=40.00n
XX1 ZN A net9 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX0 net9 B1 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX28 net9 net21 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS AOI2XB1V2_12TH40
.SUBCKT AOI2XB1V3_12TH40 A B1 B2 ZN VDD VSS
XX4 net21 B2 VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX2 ZN A VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX9 ZN B1 net25 VPW NHVT11LL_CKT W=0.71u L=40.00n
XX8 net25 net21 VSS VPW NHVT11LL_CKT W=0.71u L=40.00n
XX3 net21 B2 VDD VNW PHVT11LL_CKT W=0.26u L=40.00n
XX1 ZN A net9 VNW PHVT11LL_CKT W=0.86u L=40.00n
XX0 net9 B1 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX28 net9 net21 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
.ENDS AOI2XB1V3_12TH40
.SUBCKT AOI2XB1V4_12TH40 A B1 B2 ZN VDD VSS
XX4 net21 B2 VSS VPW NHVT11LL_CKT W=0.305u L=40.00n
XX2 ZN A VSS VPW NHVT11LL_CKT W=0.57u L=40.00n
XX9 ZN B1 net25 VPW NHVT11LL_CKT W=1.01u L=40.00n
XX8 net25 net21 VSS VPW NHVT11LL_CKT W=1.01u L=40.00n
XX3 net21 B2 VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX1 ZN A net9 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 net9 B1 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX28 net9 net21 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS AOI2XB1V4_12TH40
.SUBCKT AOI2XB1V6_12TH40 A B1 B2 ZN VDD VSS
XX4 net21 B2 VSS VPW NHVT11LL_CKT W=0.44u L=40.00n
XX2 ZN A VSS VPW NHVT11LL_CKT W=0.855u L=40.00n
XX9 ZN B1 net25 VPW NHVT11LL_CKT W=1.515u L=40.00n
XX8 net25 net21 VSS VPW NHVT11LL_CKT W=1.515u L=40.00n
XX3 net21 B2 VDD VNW PHVT11LL_CKT W=0.505u L=40.00n
XX1 ZN A net9 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX0 net9 B1 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX28 net9 net21 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS AOI2XB1V6_12TH40
.SUBCKT AOI2XB1V8_12TH40 A B1 B2 ZN VDD VSS
XX4 net21 B2 VSS VPW NHVT11LL_CKT W=0.59u L=40.00n
XX2 ZN A VSS VPW NHVT11LL_CKT W=1.14u L=40.00n
XX9 ZN B1 net25 VPW NHVT11LL_CKT W=2.02u L=40.00n
XX8 net25 net21 VSS VPW NHVT11LL_CKT W=2.02u L=40.00n
XX3 net21 B2 VDD VNW PHVT11LL_CKT W=0.67u L=40.00n
XX1 ZN A net9 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX0 net9 B1 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX28 net9 net21 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS AOI2XB1V8_12TH40
.SUBCKT AOI31V0_12TH40 A1 A2 A3 B ZN VDD VSS
XX3 net22 A3 VSS VPW NHVT11LL_CKT W=0.305u L=40.00n
XX2 ZN B VSS VPW NHVT11LL_CKT W=0.125u L=40.00n
XX9 ZN A1 net34 VPW NHVT11LL_CKT W=0.305u L=40.00n
XX8 net34 A2 net22 VPW NHVT11LL_CKT W=0.305u L=40.00n
XX4 net6 A3 VDD VNW PHVT11LL_CKT W=0.265u L=40.00n
XX1 ZN B net6 VNW PHVT11LL_CKT W=0.265u L=40.00n
XX0 net6 A2 VDD VNW PHVT11LL_CKT W=0.265u L=40.00n
XX28 net6 A1 VDD VNW PHVT11LL_CKT W=0.265u L=40.00n
.ENDS AOI31V0_12TH40
.SUBCKT AOI31V12_12TH40 A1 A2 A3 B ZN VDD VSS
XX3 net22 A3 VSS VPW NHVT11LL_CKT W=3.66u L=40.00n
XX2 ZN B VSS VPW NHVT11LL_CKT W=1.5u L=40.00n
XX9 ZN A1 net34 VPW NHVT11LL_CKT W=3.66u L=40.00n
XX8 net34 A2 net22 VPW NHVT11LL_CKT W=3.66u L=40.00n
XX4 net6 A3 VDD VNW PHVT11LL_CKT W=3.21u L=40.00n
XX1 ZN B net6 VNW PHVT11LL_CKT W=3.21u L=40.00n
XX0 net6 A2 VDD VNW PHVT11LL_CKT W=3.21u L=40.00n
XX28 net6 A1 VDD VNW PHVT11LL_CKT W=3.21u L=40.00n
.ENDS AOI31V12_12TH40
.SUBCKT AOI31V1_12TH40 A1 A2 A3 B ZN VDD VSS
XX3 net22 A3 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX2 ZN B VSS VPW NHVT11LL_CKT W=0.175u L=40.00n
XX9 ZN A1 net34 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX8 net34 A2 net22 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX4 net6 A3 VDD VNW PHVT11LL_CKT W=0.375u L=40.00n
XX1 ZN B net6 VNW PHVT11LL_CKT W=0.375u L=40.00n
XX0 net6 A2 VDD VNW PHVT11LL_CKT W=0.375u L=40.00n
XX28 net6 A1 VDD VNW PHVT11LL_CKT W=0.375u L=40.00n
.ENDS AOI31V1_12TH40
.SUBCKT AOI31V2_12TH40 A1 A2 A3 B ZN VDD VSS
XX3 net22 A3 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX2 ZN B VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX9 ZN A1 net34 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX8 net34 A2 net22 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX4 net6 A3 VDD VNW PHVT11LL_CKT W=535.00n L=40.00n
XX1 ZN B net6 VNW PHVT11LL_CKT W=535.00n L=40.00n
XX0 net6 A2 VDD VNW PHVT11LL_CKT W=535.00n L=40.00n
XX28 net6 A1 VDD VNW PHVT11LL_CKT W=535.00n L=40.00n
.ENDS AOI31V2_12TH40
.SUBCKT AOI31V3_12TH40 A1 A2 A3 B ZN VDD VSS
XX3 net22 A3 VSS VPW NHVT11LL_CKT W=0.86u L=40.00n
XX2 ZN B VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX9 ZN A1 net34 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX8 net34 A2 net22 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX4 net6 A3 VDD VNW PHVT11LL_CKT W=0.75u L=40.00n
XX1 ZN B net6 VNW PHVT11LL_CKT W=0.75u L=40.00n
XX0 net6 A2 VDD VNW PHVT11LL_CKT W=0.75u L=40.00n
XX28 net6 A1 VDD VNW PHVT11LL_CKT W=0.75u L=40.00n
.ENDS AOI31V3_12TH40
.SUBCKT AOI31V4_12TH40 A1 A2 A3 B ZN VDD VSS
XX3 net22 A3 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX2 ZN B VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX9 ZN A1 net34 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX8 net34 A2 net22 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX4 net6 A3 VDD VNW PHVT11LL_CKT W=1.07u L=40.00n
XX1 ZN B net6 VNW PHVT11LL_CKT W=1.07u L=40.00n
XX0 net6 A2 VDD VNW PHVT11LL_CKT W=1.07u L=40.00n
XX28 net6 A1 VDD VNW PHVT11LL_CKT W=1.07u L=40.00n
.ENDS AOI31V4_12TH40
.SUBCKT AOI31V6_12TH40 A1 A2 A3 B ZN VDD VSS
XX3 net22 A3 VSS VPW NHVT11LL_CKT W=1.83u L=40.00n
XX2 ZN B VSS VPW NHVT11LL_CKT W=0.75u L=40.00n
XX9 ZN A1 net34 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX8 net34 A2 net22 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX4 net6 A3 VDD VNW PHVT11LL_CKT W=1.605u L=40.00n
XX1 ZN B net6 VNW PHVT11LL_CKT W=1.605u L=40.00n
XX0 net6 A2 VDD VNW PHVT11LL_CKT W=1.605u L=40.00n
XX28 net6 A1 VDD VNW PHVT11LL_CKT W=1.605u L=40.00n
.ENDS AOI31V6_12TH40
.SUBCKT AOI31V8_12TH40 A1 A2 A3 B ZN VDD VSS
XX3 net22 A3 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX2 ZN B VSS VPW NHVT11LL_CKT W=1u L=40.00n
XX9 ZN A1 net34 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX8 net34 A2 net22 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX4 net6 A3 VDD VNW PHVT11LL_CKT W=2.14u L=40.00n
XX1 ZN B net6 VNW PHVT11LL_CKT W=2.14u L=40.00n
XX0 net6 A2 VDD VNW PHVT11LL_CKT W=2.14u L=40.00n
XX28 net6 A1 VDD VNW PHVT11LL_CKT W=2.14u L=40.00n
.ENDS AOI31V8_12TH40
.SUBCKT AOI32V0_12TH40 A1 A2 A3 B1 B2 ZN VDD VSS
XX5 net056 B2 VSS VPW NHVT11LL_CKT W=0.22u L=40.00n
XX8 net6 A2 net18 VPW NHVT11LL_CKT W=0.305u L=40.00n
XX9 ZN A1 net6 VPW NHVT11LL_CKT W=0.305u L=40.00n
XX2 ZN B1 net056 VPW NHVT11LL_CKT W=0.22u L=40.00n
XX3 net18 A3 VSS VPW NHVT11LL_CKT W=0.305u L=40.00n
XX6 ZN B1 net34 VNW PHVT11LL_CKT W=0.265u L=40.00n
XX1 ZN B2 net34 VNW PHVT11LL_CKT W=0.265u L=40.00n
XX0 net34 A2 VDD VNW PHVT11LL_CKT W=0.265u L=40.00n
XX4 net34 A3 VDD VNW PHVT11LL_CKT W=0.265u L=40.00n
XX28 net34 A1 VDD VNW PHVT11LL_CKT W=0.265u L=40.00n
.ENDS AOI32V0_12TH40
.SUBCKT AOI32V12_12TH40 A1 A2 A3 B1 B2 ZN VDD VSS
XX5 net056 B2 VSS VPW NHVT11LL_CKT W=2.64u L=40.00n
XX8 net6 A2 net18 VPW NHVT11LL_CKT W=3.66u L=40.00n
XX9 ZN A1 net6 VPW NHVT11LL_CKT W=3.66u L=40.00n
XX2 ZN B1 net056 VPW NHVT11LL_CKT W=2.64u L=40.00n
XX3 net18 A3 VSS VPW NHVT11LL_CKT W=3.66u L=40.00n
XX6 ZN B1 net34 VNW PHVT11LL_CKT W=3.21u L=40.00n
XX1 ZN B2 net34 VNW PHVT11LL_CKT W=3.21u L=40.00n
XX0 net34 A2 VDD VNW PHVT11LL_CKT W=3.21u L=40.00n
XX4 net34 A3 VDD VNW PHVT11LL_CKT W=3.21u L=40.00n
XX28 net34 A1 VDD VNW PHVT11LL_CKT W=3.21u L=40.00n
.ENDS AOI32V12_12TH40
.SUBCKT AOI32V1_12TH40 A1 A2 A3 B1 B2 ZN VDD VSS
XX5 net056 B2 VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX8 net6 A2 net18 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX9 ZN A1 net6 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX2 ZN B1 net056 VPW NHVT11LL_CKT W=0.31u L=40.00n
XX3 net18 A3 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX6 ZN B1 net34 VNW PHVT11LL_CKT W=0.375u L=40.00n
XX1 ZN B2 net34 VNW PHVT11LL_CKT W=0.375u L=40.00n
XX0 net34 A2 VDD VNW PHVT11LL_CKT W=0.375u L=40.00n
XX4 net34 A3 VDD VNW PHVT11LL_CKT W=0.375u L=40.00n
XX28 net34 A1 VDD VNW PHVT11LL_CKT W=0.375u L=40.00n
.ENDS AOI32V1_12TH40
.SUBCKT AOI32V2_12TH40 A1 A2 A3 B1 B2 ZN VDD VSS
XX5 net056 B2 VSS VPW NHVT11LL_CKT W=440.00n L=40.00n
XX8 net6 A2 net18 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX9 ZN A1 net6 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX2 ZN B1 net056 VPW NHVT11LL_CKT W=440.00n L=40.00n
XX3 net18 A3 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX6 ZN B1 net34 VNW PHVT11LL_CKT W=535.00n L=40.00n
XX1 ZN B2 net34 VNW PHVT11LL_CKT W=535.00n L=40.00n
XX0 net34 A2 VDD VNW PHVT11LL_CKT W=535.00n L=40.00n
XX4 net34 A3 VDD VNW PHVT11LL_CKT W=535.00n L=40.00n
XX28 net34 A1 VDD VNW PHVT11LL_CKT W=535.00n L=40.00n
.ENDS AOI32V2_12TH40
.SUBCKT AOI32V3_12TH40 A1 A2 A3 B1 B2 ZN VDD VSS
XX5 net056 B2 VSS VPW NHVT11LL_CKT W=0.62u L=40.00n
XX8 net6 A2 net18 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX9 ZN A1 net6 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX2 ZN B1 net056 VPW NHVT11LL_CKT W=0.62u L=40.00n
XX3 net18 A3 VSS VPW NHVT11LL_CKT W=0.86u L=40.00n
XX6 ZN B1 net34 VNW PHVT11LL_CKT W=0.75u L=40.00n
XX1 ZN B2 net34 VNW PHVT11LL_CKT W=0.75u L=40.00n
XX0 net34 A2 VDD VNW PHVT11LL_CKT W=0.75u L=40.00n
XX4 net34 A3 VDD VNW PHVT11LL_CKT W=0.75u L=40.00n
XX28 net34 A1 VDD VNW PHVT11LL_CKT W=0.75u L=40.00n
.ENDS AOI32V3_12TH40
.SUBCKT AOI32V4_12TH40 A1 A2 A3 B1 B2 ZN VDD VSS
XX5 net056 B2 VSS VPW NHVT11LL_CKT W=0.88u L=40.00n
XX8 net6 A2 net18 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX9 ZN A1 net6 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX2 ZN B1 net056 VPW NHVT11LL_CKT W=0.88u L=40.00n
XX3 net18 A3 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX6 ZN B1 net34 VNW PHVT11LL_CKT W=1.07u L=40.00n
XX1 ZN B2 net34 VNW PHVT11LL_CKT W=1.07u L=40.00n
XX0 net34 A2 VDD VNW PHVT11LL_CKT W=1.07u L=40.00n
XX4 net34 A3 VDD VNW PHVT11LL_CKT W=1.07u L=40.00n
XX28 net34 A1 VDD VNW PHVT11LL_CKT W=1.07u L=40.00n
.ENDS AOI32V4_12TH40
.SUBCKT AOI32V6_12TH40 A1 A2 A3 B1 B2 ZN VDD VSS
XX5 net056 B2 VSS VPW NHVT11LL_CKT W=1.32u L=40.00n
XX8 net6 A2 net18 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX9 ZN A1 net6 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX2 ZN B1 net056 VPW NHVT11LL_CKT W=1.32u L=40.00n
XX3 net18 A3 VSS VPW NHVT11LL_CKT W=1.83u L=40.00n
XX6 ZN B1 net34 VNW PHVT11LL_CKT W=1.605u L=40.00n
XX1 ZN B2 net34 VNW PHVT11LL_CKT W=1.605u L=40.00n
XX0 net34 A2 VDD VNW PHVT11LL_CKT W=1.605u L=40.00n
XX4 net34 A3 VDD VNW PHVT11LL_CKT W=1.605u L=40.00n
XX28 net34 A1 VDD VNW PHVT11LL_CKT W=1.605u L=40.00n
.ENDS AOI32V6_12TH40
.SUBCKT AOI32V8_12TH40 A1 A2 A3 B1 B2 ZN VDD VSS
XX5 net056 B2 VSS VPW NHVT11LL_CKT W=1.76u L=40.00n
XX8 net6 A2 net18 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX9 ZN A1 net6 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX2 ZN B1 net056 VPW NHVT11LL_CKT W=1.76u L=40.00n
XX3 net18 A3 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX6 ZN B1 net34 VNW PHVT11LL_CKT W=2.14u L=40.00n
XX1 ZN B2 net34 VNW PHVT11LL_CKT W=2.14u L=40.00n
XX0 net34 A2 VDD VNW PHVT11LL_CKT W=2.14u L=40.00n
XX4 net34 A3 VDD VNW PHVT11LL_CKT W=2.14u L=40.00n
XX28 net34 A1 VDD VNW PHVT11LL_CKT W=2.14u L=40.00n
.ENDS AOI32V8_12TH40
.SUBCKT AOI33V1_12TH40 A1 A2 A3 B1 B2 B3 ZN VDD VSS
XX11 net028 B3 VSS VPW NHVT11LL_CKT W=430.00n L=40.00n
XX5 net056 B2 net028 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX8 net6 A2 net18 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX9 ZN A1 net6 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX2 ZN B1 net056 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX3 net18 A3 VSS VPW NHVT11LL_CKT W=430.00n L=40.00n
XX12 ZN B3 net34 VNW PHVT11LL_CKT W=380.00n L=40.00n
XX6 ZN B1 net34 VNW PHVT11LL_CKT W=380.00n L=40.00n
XX1 ZN B2 net34 VNW PHVT11LL_CKT W=380.00n L=40.00n
XX0 net34 A2 VDD VNW PHVT11LL_CKT W=380.00n L=40.00n
XX4 net34 A3 VDD VNW PHVT11LL_CKT W=380.00n L=40.00n
XX28 net34 A1 VDD VNW PHVT11LL_CKT W=380.00n L=40.00n
.ENDS AOI33V1_12TH40
.SUBCKT AOI33V2_12TH40 A1 A2 A3 B1 B2 B3 ZN VDD VSS
XX0 net43 A2 VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX4 net43 A3 VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX28 net43 A1 VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX12 ZN B3 net43 VNW PHVT11LL_CKT W=540.00n L=40.00n
XX6 ZN B1 net43 VNW PHVT11LL_CKT W=540.00n L=40.00n
XX1 ZN B2 net43 VNW PHVT11LL_CKT W=540.00n L=40.00n
XX3 net52 A3 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX11 net72 B3 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX5 net68 B2 net72 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX8 net64 A2 net52 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX9 ZN A1 net64 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX2 ZN B1 net68 VPW NHVT11LL_CKT W=610.00n L=40.00n
.ENDS AOI33V2_12TH40
.SUBCKT AOI33V4_12TH40 A1 A2 A3 B1 B2 B3 ZN VDD VSS
XX0 net43 A2 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX4 net43 A3 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX28 net43 A1 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX12 ZN B3 net43 VNW PHVT11LL_CKT W=1.08u L=40.00n
XX6 ZN B1 net43 VNW PHVT11LL_CKT W=1.08u L=40.00n
XX1 ZN B2 net43 VNW PHVT11LL_CKT W=1.08u L=40.00n
XX3 net52 A3 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX11 net72 B3 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX5 net68 B2 net72 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX8 net64 A2 net52 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX9 ZN A1 net64 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX2 ZN B1 net68 VPW NHVT11LL_CKT W=1.22u L=40.00n
.ENDS AOI33V4_12TH40
.SUBCKT AOI33V8_12TH40 A1 A2 A3 B1 B2 B3 ZN VDD VSS
XX0 net43 A2 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
XX4 net43 A3 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
XX28 net43 A1 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
XX12 ZN B3 net43 VNW PHVT11LL_CKT W=2.16u L=40.00n
XX6 ZN B1 net43 VNW PHVT11LL_CKT W=2.16u L=40.00n
XX1 ZN B2 net43 VNW PHVT11LL_CKT W=2.16u L=40.00n
XX3 net52 A3 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX11 net72 B3 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX5 net68 B2 net72 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX8 net64 A2 net52 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX9 ZN A1 net64 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX2 ZN B1 net68 VPW NHVT11LL_CKT W=2.44u L=40.00n
.ENDS AOI33V8_12TH40
.SUBCKT BENCV12_12TH40 A MI0 MI1 MI2 S X2 VDD VSS
XX17 A net_413 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX16 net_413 net_349 VDD VNW PHVT11LL_CKT W=0.91u L=40.00n
XX15 net_349 MI0 net_352 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX14 net_349 net100 VDD VNW PHVT11LL_CKT W=0.26u L=40.00n
XX13 net_352 MI1 VDD VNW PHVT11LL_CKT W=0.48u L=40.00n
XX11 net106 net108 net_412 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX9 X2 net_401 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX8 net_401 net_412 VDD VNW PHVT11LL_CKT W=0.91u L=40.00n
XX10 net110 MI1 net_412 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX5 net_377 net_313 VDD VNW PHVT11LL_CKT W=0.91u L=40.00n
XX6 S net_377 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX4 net_313 net110 net_316 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX3 net_313 MI2 VDD VNW PHVT11LL_CKT W=0.26u L=40.00n
XX2 net_316 net108 VDD VNW PHVT11LL_CKT W=0.48u L=40.00n
XX0 net110 MI0 VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
XX7 net108 MI1 VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX1 net106 net110 VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
XX12 net100 MI2 VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX22 net_425 MI0 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX20 net_349 net100 net_425 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX18 A net_413 VSS VPW NHVT11LL_CKT W=3.21u L=40.00n
XX19 net_413 net_349 VSS VPW NHVT11LL_CKT W=0.8u L=40.00n
XX28 net106 MI1 net_412 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX25 X2 net_401 VSS VPW NHVT11LL_CKT W=3.21u L=40.00n
XX26 net_401 net_412 VSS VPW NHVT11LL_CKT W=0.8u L=40.00n
XX27 net110 net108 net_412 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX35 net_389 net110 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX34 net_389 net108 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX33 net_313 MI2 net_389 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX36 S net_377 VSS VPW NHVT11LL_CKT W=3.21u L=40.00n
XX31 net_377 net_313 VSS VPW NHVT11LL_CKT W=0.8u L=40.00n
XX30 net106 net110 VSS VPW NHVT11LL_CKT W=410.00n L=40.00n
XX29 net110 MI0 VSS VPW NHVT11LL_CKT W=410.00n L=40.00n
XX21 net_425 MI1 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX24 net108 MI1 VSS VPW NHVT11LL_CKT W=0.39u L=40.00n
XX23 net100 MI2 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
.ENDS BENCV12_12TH40
.SUBCKT BENCV16_12TH40 A MI0 MI1 MI2 S X2 VDD VSS
XX17 A net_413 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX16 net_413 net_349 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX15 net_349 MI0 net_352 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX14 net_349 net100 VDD VNW PHVT11LL_CKT W=0.325u L=40.00n
XX13 net_352 MI1 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX11 net106 net108 net_412 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX9 X2 net_401 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX8 net_401 net_412 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX10 net110 MI1 net_412 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX5 net_377 net_313 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX6 S net_377 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX4 net_313 net110 net_316 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX3 net_313 MI2 VDD VNW PHVT11LL_CKT W=0.325u L=40.00n
XX2 net_316 net108 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net110 MI0 VDD VNW PHVT11LL_CKT W=0.535u L=40.00n
XX7 net108 MI1 VDD VNW PHVT11LL_CKT W=470.00n L=40.00n
XX1 net106 net110 VDD VNW PHVT11LL_CKT W=0.535u L=40.00n
XX12 net100 MI2 VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX22 net_425 MI0 VSS VPW NHVT11LL_CKT W=0.505u L=40.00n
XX20 net_349 net100 net_425 VPW NHVT11LL_CKT W=0.505u L=40.00n
XX18 A net_413 VSS VPW NHVT11LL_CKT W=4.28u L=40.00n
XX19 net_413 net_349 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX28 net106 MI1 net_412 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX25 X2 net_401 VSS VPW NHVT11LL_CKT W=4.28u L=40.00n
XX26 net_401 net_412 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX27 net110 net108 net_412 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX35 net_389 net110 VSS VPW NHVT11LL_CKT W=0.505u L=40.00n
XX34 net_389 net108 VSS VPW NHVT11LL_CKT W=0.505u L=40.00n
XX33 net_313 MI2 net_389 VPW NHVT11LL_CKT W=0.505u L=40.00n
XX36 S net_377 VSS VPW NHVT11LL_CKT W=4.28u L=40.00n
XX31 net_377 net_313 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX30 net106 net110 VSS VPW NHVT11LL_CKT W=0.44u L=40.00n
XX29 net110 MI0 VSS VPW NHVT11LL_CKT W=0.44u L=40.00n
XX21 net_425 MI1 VSS VPW NHVT11LL_CKT W=0.505u L=40.00n
XX24 net108 MI1 VSS VPW NHVT11LL_CKT W=410.00n L=40.00n
XX23 net100 MI2 VSS VPW NHVT11LL_CKT W=140.00n L=40.00n
.ENDS BENCV16_12TH40
.SUBCKT BENCV20_12TH40 A MI0 MI1 MI2 S X2 VDD VSS
XX17 A net_413 VDD VNW PHVT11LL_CKT W=6.1u L=40.00n
XX16 net_413 net_349 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX15 net_349 MI0 net_352 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX14 net_349 net100 VDD VNW PHVT11LL_CKT W=0.325u L=40.00n
XX13 net_352 MI1 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX11 net106 net108 net_412 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX9 X2 net_401 VDD VNW PHVT11LL_CKT W=6.1u L=40.00n
XX8 net_401 net_412 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX10 net110 MI1 net_412 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX5 net_377 net_313 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX6 S net_377 VDD VNW PHVT11LL_CKT W=6.1u L=40.00n
XX4 net_313 net110 net_316 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX3 net_313 MI2 VDD VNW PHVT11LL_CKT W=0.325u L=40.00n
XX2 net_316 net108 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net110 MI0 VDD VNW PHVT11LL_CKT W=0.58u L=40.00n
XX7 net108 MI1 VDD VNW PHVT11LL_CKT W=470.00n L=40.00n
XX1 net106 net110 VDD VNW PHVT11LL_CKT W=0.58u L=40.00n
XX12 net100 MI2 VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX22 net_425 MI0 VSS VPW NHVT11LL_CKT W=0.505u L=40.00n
XX20 net_349 net100 net_425 VPW NHVT11LL_CKT W=0.505u L=40.00n
XX18 A net_413 VSS VPW NHVT11LL_CKT W=5.35u L=40.00n
XX19 net_413 net_349 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX28 net106 MI1 net_412 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX25 X2 net_401 VSS VPW NHVT11LL_CKT W=5.35u L=40.00n
XX26 net_401 net_412 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX27 net110 net108 net_412 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX35 net_389 net110 VSS VPW NHVT11LL_CKT W=0.505u L=40.00n
XX34 net_389 net108 VSS VPW NHVT11LL_CKT W=0.505u L=40.00n
XX33 net_313 MI2 net_389 VPW NHVT11LL_CKT W=0.505u L=40.00n
XX36 S net_377 VSS VPW NHVT11LL_CKT W=5.35u L=40.00n
XX31 net_377 net_313 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX30 net106 net110 VSS VPW NHVT11LL_CKT W=0.48u L=40.00n
XX29 net110 MI0 VSS VPW NHVT11LL_CKT W=0.48u L=40.00n
XX21 net_425 MI1 VSS VPW NHVT11LL_CKT W=0.505u L=40.00n
XX24 net108 MI1 VSS VPW NHVT11LL_CKT W=410.00n L=40.00n
XX23 net100 MI2 VSS VPW NHVT11LL_CKT W=140.00n L=40.00n
.ENDS BENCV20_12TH40
.SUBCKT BENCV32_12TH40 A MI0 MI1 MI2 S X2 VDD VSS
XX17 A net_413 VDD VNW PHVT11LL_CKT W=9.76u L=40.00n
XX16 net_413 net_349 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX15 net_349 MI0 net_352 VNW PHVT11LL_CKT W=0.9u L=40.00n
XX14 net_349 net100 VDD VNW PHVT11LL_CKT W=0.47u L=40.00n
XX13 net_352 MI1 VDD VNW PHVT11LL_CKT W=0.9u L=40.00n
XX11 net106 net108 net_412 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX9 X2 net_401 VDD VNW PHVT11LL_CKT W=9.76u L=40.00n
XX8 net_401 net_412 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX10 net110 MI1 net_412 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX5 net_377 net_313 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX6 S net_377 VDD VNW PHVT11LL_CKT W=9.76u L=40.00n
XX4 net_313 net110 net_316 VNW PHVT11LL_CKT W=0.9u L=40.00n
XX3 net_313 MI2 VDD VNW PHVT11LL_CKT W=0.47u L=40.00n
XX2 net_316 net108 VDD VNW PHVT11LL_CKT W=0.9u L=40.00n
XX0 net110 MI0 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX7 net108 MI1 VDD VNW PHVT11LL_CKT W=0.57u L=40.00n
XX1 net106 net110 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX12 net100 MI2 VDD VNW PHVT11LL_CKT W=0.34u L=40.00n
XX22 net_425 MI0 VSS VPW NHVT11LL_CKT W=0.74u L=40.00n
XX20 net_349 net100 net_425 VPW NHVT11LL_CKT W=0.74u L=40.00n
XX18 A net_413 VSS VPW NHVT11LL_CKT W=8.56u L=40.00n
XX19 net_413 net_349 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX28 net106 MI1 net_412 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX25 X2 net_401 VSS VPW NHVT11LL_CKT W=8.56u L=40.00n
XX26 net_401 net_412 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX27 net110 net108 net_412 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX35 net_389 net110 VSS VPW NHVT11LL_CKT W=0.74u L=40.00n
XX34 net_389 net108 VSS VPW NHVT11LL_CKT W=0.74u L=40.00n
XX33 net_313 MI2 net_389 VPW NHVT11LL_CKT W=0.74u L=40.00n
XX36 S net_377 VSS VPW NHVT11LL_CKT W=8.56u L=40.00n
XX31 net_377 net_313 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX30 net106 net110 VSS VPW NHVT11LL_CKT W=0.505u L=40.00n
XX29 net110 MI0 VSS VPW NHVT11LL_CKT W=0.505u L=40.00n
XX21 net_425 MI1 VSS VPW NHVT11LL_CKT W=0.74u L=40.00n
XX24 net108 MI1 VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX23 net100 MI2 VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
.ENDS BENCV32_12TH40
.SUBCKT BENCV4_12TH40 A MI0 MI1 MI2 S X2 VDD VSS
XX33 net_67 MI0 net_119 VPW NHVT11LL_CKT W=505.00n L=40.00n
XX30 net106 net110 VSS VPW NHVT11LL_CKT W=410.00n L=40.00n
XX29 net110 MI0 VSS VPW NHVT11LL_CKT W=410.00n L=40.00n
XX28 net106 net108 net_82 VPW NHVT11LL_CKT W=410.00n L=40.00n
XX27 net110 MI1 net_82 VPW NHVT11LL_CKT W=410.00n L=40.00n
XX25 X2 net_82 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX24 net108 MI1 VSS VPW NHVT11LL_CKT W=410.00n L=40.00n
XX23 net100 MI2 VSS VPW NHVT11LL_CKT W=140.00n L=40.00n
XX37 net_107 MI2 VSS VPW NHVT11LL_CKT W=285.00n L=40.00n
XX38 net_103 net108 VSS VPW NHVT11LL_CKT W=505.00n L=40.00n
XX39 net_107 net110 net_103 VPW NHVT11LL_CKT W=505.00n L=40.00n
XX18 A net_107 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX36 S net_67 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX34 net_119 MI1 VSS VPW NHVT11LL_CKT W=505.00n L=40.00n
XX35 net_67 net100 VSS VPW NHVT11LL_CKT W=285.00n L=40.00n
XX10 net110 net108 net_82 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX0 net110 MI0 VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
XX4 net_67 net100 net_18 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX2 net_18 MI0 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX3 net_18 MI1 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX11 net106 MI1 net_82 VNW PHVT11LL_CKT W=500.00n L=40.00n
XX7 net108 MI1 VDD VNW PHVT11LL_CKT W=470.00n L=40.00n
XX19 net_62 net108 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 net106 net110 VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
XX6 S net_67 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX17 A net_107 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX9 X2 net_82 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX20 net_62 net110 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX21 net_107 MI2 net_62 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX12 net100 MI2 VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
.ENDS BENCV4_12TH40
.SUBCKT BENCV6_12TH40 A MI0 MI1 MI2 S X2 VDD VSS
XX18 A net_163 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX20 net_179 net100 net_151 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX19 net_163 net_179 VSS VPW NHVT11LL_CKT W=0.45u L=40.00n
XX21 net_151 MI1 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX22 net_151 MI0 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX25 X2 net_143 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX26 net_143 net_138 VSS VPW NHVT11LL_CKT W=0.45u L=40.00n
XX27 net110 net108 net_138 VPW NHVT11LL_CKT W=0.27u L=40.00n
XX28 net106 MI1 net_138 VPW NHVT11LL_CKT W=0.27u L=40.00n
XX31 net_131 net_219 VSS VPW NHVT11LL_CKT W=0.45u L=40.00n
XX33 net_219 MI2 net_123 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX34 net_123 net108 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX35 net_123 net110 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX36 S net_131 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX30 net106 net110 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX29 net110 MI0 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX24 net108 MI1 VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX23 net100 MI2 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX13 net_182 MI1 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX14 net_179 net100 VDD VNW PHVT11LL_CKT W=0.165u L=40.00n
XX15 net_179 MI0 net_182 VNW PHVT11LL_CKT W=0.305u L=40.00n
XX16 net_163 net_179 VDD VNW PHVT11LL_CKT W=0.515u L=40.00n
XX17 A net_163 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX3 net_219 MI2 VDD VNW PHVT11LL_CKT W=0.165u L=40.00n
XX2 net_222 net108 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX11 net106 net108 net_138 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX5 net_131 net_219 VDD VNW PHVT11LL_CKT W=0.515u L=40.00n
XX9 X2 net_143 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX6 S net_131 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX10 net110 MI1 net_138 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX4 net_219 net110 net_222 VNW PHVT11LL_CKT W=0.305u L=40.00n
XX8 net_143 net_138 VDD VNW PHVT11LL_CKT W=0.515u L=40.00n
XX0 net110 MI0 VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX7 net108 MI1 VDD VNW PHVT11LL_CKT W=0.32u L=40.00n
XX1 net106 net110 VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX12 net100 MI2 VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
.ENDS BENCV6_12TH40
.SUBCKT BENCV8_12TH40 A MI0 MI1 MI2 S X2 VDD VSS
XX17 A net_413 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX16 net_413 net_349 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX15 net_349 MI0 net_352 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX14 net_349 net100 VDD VNW PHVT11LL_CKT W=0.18u L=40.00n
XX13 net_352 MI1 VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX11 net106 net108 net_412 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX9 X2 net_401 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX8 net_401 net_412 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX10 net110 MI1 net_412 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX5 net_377 net_313 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX6 S net_377 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX4 net_313 net110 net_316 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX3 net_313 MI2 VDD VNW PHVT11LL_CKT W=0.18u L=40.00n
XX2 net_316 net108 VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX0 net110 MI0 VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX7 net108 MI1 VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX1 net106 net110 VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX12 net100 MI2 VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX22 net_425 MI0 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX20 net_349 net100 net_425 VPW NHVT11LL_CKT W=0.27u L=40.00n
XX18 A net_413 VSS VPW NHVT11LL_CKT W=2.14u L=40.00n
XX19 net_413 net_349 VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX28 net106 MI1 net_412 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX25 X2 net_401 VSS VPW NHVT11LL_CKT W=2.14u L=40.00n
XX26 net_401 net_412 VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX27 net110 net108 net_412 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX35 net_389 net110 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX34 net_389 net108 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX33 net_313 MI2 net_389 VPW NHVT11LL_CKT W=0.27u L=40.00n
XX36 S net_377 VSS VPW NHVT11LL_CKT W=2.14u L=40.00n
XX31 net_377 net_313 VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX30 net106 net110 VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX29 net110 MI0 VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX21 net_425 MI1 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX24 net108 MI1 VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX23 net100 MI2 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
.ENDS BENCV8_12TH40
.SUBCKT BMUXNV1_12TH40 A MI0 MI1 PPN S X2 VDD VSS
XX23 PPN net076 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX21 X2N X2 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX19 MSAD0 X2 net076 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX18 MASD1 X2N net076 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX15 SN MI0N MSAD0 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX14 AN MI0 MSAD0 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX9 SN MI1N MASD1 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX8 AN MI1 MASD1 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX4 MI1N MI1 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX3 MI0N MI0 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX2 SN S VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX7 AN A VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX20 X2N X2 VDD VNW PHVT11LL_CKT W=0.28u L=40.00n
XX22 PPN net076 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX17 MSAD0 X2N net076 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX16 MASD1 X2 net076 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX11 SN MI1 MASD1 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX10 AN MI1N MASD1 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX13 SN MI0 MSAD0 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX5 MI1N MI1 VDD VNW PHVT11LL_CKT W=0.28u L=40.00n
XX0 MI0N MI0 VDD VNW PHVT11LL_CKT W=0.28u L=40.00n
XX12 AN MI0N MSAD0 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX1 SN S VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX6 AN A VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
.ENDS BMUXNV1_12TH40
.SUBCKT BMUXNV2_12TH40 A MI0 MI1 PPN S X2 VDD VSS
XX23 PPN net076 VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX21 X2N X2 VSS VPW NHVT11LL_CKT W=285.00n L=40.00n
XX19 MSAD0 X2 net076 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX18 MASD1 X2N net076 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX15 SN MI0N MSAD0 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX14 AN MI0 MSAD0 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX9 SN MI1N MASD1 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX8 AN MI1 MASD1 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX4 MI1N MI1 VSS VPW NHVT11LL_CKT W=285.00n L=40.00n
XX3 MI0N MI0 VSS VPW NHVT11LL_CKT W=285.00n L=40.00n
XX2 SN S VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX7 AN A VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX20 X2N X2 VDD VNW PHVT11LL_CKT W=325.00n L=40.00n
XX22 PPN net076 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX17 MSAD0 X2N net076 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX16 MASD1 X2 net076 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX11 SN MI1 MASD1 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX10 AN MI1N MASD1 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX13 SN MI0 MSAD0 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX5 MI1N MI1 VDD VNW PHVT11LL_CKT W=325.00n L=40.00n
XX0 MI0N MI0 VDD VNW PHVT11LL_CKT W=325.00n L=40.00n
XX12 AN MI0N MSAD0 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX1 SN S VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX6 AN A VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
.ENDS BMUXNV2_12TH40
.SUBCKT BMUXNV3_12TH40 A MI0 MI1 PPN S X2 VDD VSS
XX23 PPN net076 VSS VPW NHVT11LL_CKT W=0.76u L=40.00n
XX21 X2N X2 VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX19 MSAD0 X2 net076 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX18 MASD1 X2N net076 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX15 SN MI0N MSAD0 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX14 AN MI0 MSAD0 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX9 SN MI1N MASD1 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX8 AN MI1 MASD1 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX4 MI1N MI1 VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX3 MI0N MI0 VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX2 SN S VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX7 AN A VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX20 X2N X2 VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX22 PPN net076 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX17 MSAD0 X2N net076 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX16 MASD1 X2 net076 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX11 SN MI1 MASD1 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX10 AN MI1N MASD1 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX13 SN MI0 MSAD0 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX5 MI1N MI1 VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX0 MI0N MI0 VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX12 AN MI0N MSAD0 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX1 SN S VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX6 AN A VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
.ENDS BMUXNV3_12TH40
.SUBCKT BMUXNV4_12TH40 A MI0 MI1 PPN S X2 VDD VSS
XX23 PPN net076 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX21 X2N X2 VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX19 MSAD0 X2 net076 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX18 MASD1 X2N net076 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX15 SN MI0N MSAD0 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX14 AN MI0 MSAD0 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX9 SN MI1N MASD1 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX8 AN MI1 MASD1 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX4 MI1N MI1 VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX3 MI0N MI0 VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX2 SN S VSS VPW NHVT11LL_CKT W=0.46u L=40.00n
XX7 AN A VSS VPW NHVT11LL_CKT W=0.46u L=40.00n
XX20 X2N X2 VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX22 PPN net076 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX17 MSAD0 X2N net076 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX16 MASD1 X2 net076 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX11 SN MI1 MASD1 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX10 AN MI1N MASD1 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX13 SN MI0 MSAD0 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX5 MI1N MI1 VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX0 MI0N MI0 VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX12 AN MI0N MSAD0 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX1 SN S VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX6 AN A VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
.ENDS BMUXNV4_12TH40
.SUBCKT BMUXV1_12TH40 A MI0 MI1 PP S X2 VDD VSS
XX26 MASD1N MASD1 VSS VPW NHVT11LL_CKT W=0.24u L=40.00n
XX24 MSAD0N MSAD0 VSS VPW NHVT11LL_CKT W=0.24u L=40.00n
XX7 AN A VSS VPW NHVT11LL_CKT W=0.24u L=40.00n
XX2 SN S VSS VPW NHVT11LL_CKT W=0.24u L=40.00n
XX3 MI0N MI0 VSS VPW NHVT11LL_CKT W=0.22u L=40.00n
XX4 MI1N MI1 VSS VPW NHVT11LL_CKT W=0.22u L=40.00n
XX8 AN MI1 MASD1 VPW NHVT11LL_CKT W=0.24u L=40.00n
XX9 SN MI1N MASD1 VPW NHVT11LL_CKT W=0.24u L=40.00n
XX14 AN MI0 MSAD0 VPW NHVT11LL_CKT W=0.24u L=40.00n
XX15 SN MI0N MSAD0 VPW NHVT11LL_CKT W=0.24u L=40.00n
XX18 MASD1N X2N net54 VPW NHVT11LL_CKT W=0.24u L=40.00n
XX19 MSAD0N X2 net54 VPW NHVT11LL_CKT W=0.24u L=40.00n
XX21 X2N X2 VSS VPW NHVT11LL_CKT W=0.22u L=40.00n
XX23 PP net54 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX27 MASD1N MASD1 VDD VNW PHVT11LL_CKT W=0.29u L=40.00n
XX25 MSAD0N MSAD0 VDD VNW PHVT11LL_CKT W=0.29u L=40.00n
XX6 AN A VDD VNW PHVT11LL_CKT W=0.29u L=40.00n
XX1 SN S VDD VNW PHVT11LL_CKT W=0.29u L=40.00n
XX12 AN MI0N MSAD0 VNW PHVT11LL_CKT W=0.29u L=40.00n
XX0 MI0N MI0 VDD VNW PHVT11LL_CKT W=0.255u L=40.00n
XX5 MI1N MI1 VDD VNW PHVT11LL_CKT W=0.255u L=40.00n
XX13 SN MI0 MSAD0 VNW PHVT11LL_CKT W=0.29u L=40.00n
XX10 AN MI1N MASD1 VNW PHVT11LL_CKT W=0.29u L=40.00n
XX11 SN MI1 MASD1 VNW PHVT11LL_CKT W=0.29u L=40.00n
XX16 MASD1N X2 net54 VNW PHVT11LL_CKT W=0.29u L=40.00n
XX17 MSAD0N X2N net54 VNW PHVT11LL_CKT W=0.29u L=40.00n
XX22 PP net54 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX20 X2N X2 VDD VNW PHVT11LL_CKT W=0.255u L=40.00n
.ENDS BMUXV1_12TH40
.SUBCKT BMUXV2_12TH40 A MI0 MI1 PP S X2 VDD VSS
XX26 MASD1N MASD1 VSS VPW NHVT11LL_CKT W=300.00n L=40.00n
XX24 MSAD0N MSAD0 VSS VPW NHVT11LL_CKT W=300.00n L=40.00n
XX7 AN A VSS VPW NHVT11LL_CKT W=300.00n L=40.00n
XX2 SN S VSS VPW NHVT11LL_CKT W=300.00n L=40.00n
XX3 MI0N MI0 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX4 MI1N MI1 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX8 AN MI1 MASD1 VPW NHVT11LL_CKT W=300.00n L=40.00n
XX9 SN MI1N MASD1 VPW NHVT11LL_CKT W=300.00n L=40.00n
XX14 AN MI0 MSAD0 VPW NHVT11LL_CKT W=300.00n L=40.00n
XX15 SN MI0N MSAD0 VPW NHVT11LL_CKT W=300.00n L=40.00n
XX18 MASD1N X2N net54 VPW NHVT11LL_CKT W=300.00n L=40.00n
XX19 MSAD0N X2 net54 VPW NHVT11LL_CKT W=300.00n L=40.00n
XX21 X2N X2 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX23 PP net54 VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX27 MASD1N MASD1 VDD VNW PHVT11LL_CKT W=360.00n L=40.00n
XX25 MSAD0N MSAD0 VDD VNW PHVT11LL_CKT W=360.00n L=40.00n
XX6 AN A VDD VNW PHVT11LL_CKT W=360.00n L=40.00n
XX1 SN S VDD VNW PHVT11LL_CKT W=360.00n L=40.00n
XX12 AN MI0N MSAD0 VNW PHVT11LL_CKT W=360.00n L=40.00n
XX0 MI0N MI0 VDD VNW PHVT11LL_CKT W=290.00n L=40.00n
XX5 MI1N MI1 VDD VNW PHVT11LL_CKT W=290.00n L=40.00n
XX13 SN MI0 MSAD0 VNW PHVT11LL_CKT W=360.00n L=40.00n
XX10 AN MI1N MASD1 VNW PHVT11LL_CKT W=360.00n L=40.00n
XX11 SN MI1 MASD1 VNW PHVT11LL_CKT W=360.00n L=40.00n
XX16 MASD1N X2 net54 VNW PHVT11LL_CKT W=360.00n L=40.00n
XX17 MSAD0N X2N net54 VNW PHVT11LL_CKT W=360.00n L=40.00n
XX22 PP net54 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX20 X2N X2 VDD VNW PHVT11LL_CKT W=290.00n L=40.00n
.ENDS BMUXV2_12TH40
.SUBCKT BMUXV3_12TH40 A MI0 MI1 PP S X2 VDD VSS
XX26 MASD1N MASD1 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX24 MSAD0N MSAD0 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX7 AN A VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX2 SN S VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX3 MI0N MI0 VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX4 MI1N MI1 VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX8 AN MI1 MASD1 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX9 SN MI1N MASD1 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX14 AN MI0 MSAD0 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX15 SN MI0N MSAD0 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX18 MASD1N X2N net54 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX19 MSAD0N X2 net54 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX21 X2N X2 VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX23 PP net54 VSS VPW NHVT11LL_CKT W=0.76u L=40.00n
XX27 MASD1N MASD1 VDD VNW PHVT11LL_CKT W=0.48u L=40.00n
XX25 MSAD0N MSAD0 VDD VNW PHVT11LL_CKT W=0.48u L=40.00n
XX6 AN A VDD VNW PHVT11LL_CKT W=0.48u L=40.00n
XX1 SN S VDD VNW PHVT11LL_CKT W=0.48u L=40.00n
XX12 AN MI0N MSAD0 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX0 MI0N MI0 VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX5 MI1N MI1 VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX13 SN MI0 MSAD0 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX10 AN MI1N MASD1 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX11 SN MI1 MASD1 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX16 MASD1N X2 net54 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX17 MSAD0N X2N net54 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX22 PP net54 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX20 X2N X2 VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
.ENDS BMUXV3_12TH40
.SUBCKT BMUXV4_12TH40 A MI0 MI1 PP S X2 VDD VSS
XX26 MASD1N MASD1 VSS VPW NHVT11LL_CKT W=0.41u L=40.00n
XX24 MSAD0N MSAD0 VSS VPW NHVT11LL_CKT W=0.41u L=40.00n
XX7 AN A VSS VPW NHVT11LL_CKT W=0.41u L=40.00n
XX2 SN S VSS VPW NHVT11LL_CKT W=0.41u L=40.00n
XX3 MI0N MI0 VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX4 MI1N MI1 VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX8 AN MI1 MASD1 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX9 SN MI1N MASD1 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX14 AN MI0 MSAD0 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX15 SN MI0N MSAD0 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX18 MASD1N X2N net54 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX19 MSAD0N X2 net54 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX21 X2N X2 VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX23 PP net54 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX27 MASD1N MASD1 VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX25 MSAD0N MSAD0 VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX6 AN A VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX1 SN S VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX12 AN MI0N MSAD0 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX0 MI0N MI0 VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX5 MI1N MI1 VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX13 SN MI0 MSAD0 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX10 AN MI1N MASD1 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX11 SN MI1 MASD1 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX16 MASD1N X2 net54 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX17 MSAD0N X2N net54 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX22 PP net54 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX20 X2N X2 VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
.ENDS BMUXV4_12TH40
.SUBCKT BUFV10RD_12TH40 I Z VDD VSS
XX1 net11 I VSS VPW NHVT11LL_CKT W=1.545u L=40.00n
XX6 Z net11 VSS VPW NHVT11LL_CKT W=2.7u L=40.00n
XX0 net11 I VDD VNW PHVT11LL_CKT W=1.77u L=40.00n
XX5 Z net11 VDD VNW PHVT11LL_CKT W=3.05u L=40.00n
.ENDS BUFV10RD_12TH40
.SUBCKT BUFV10RO_12TH40 I Z VDD VSS
XX1 net26 I VDD VNW PHVT11LL_CKT W=380.00n L=40.00n
XX3 Z net26 VDD VNW PHVT11LL_CKT W=3.05u L=40.00n
XX2 net26 I VSS VPW NHVT11LL_CKT W=340.00n L=40.00n
XX0 Z net26 VSS VPW NHVT11LL_CKT W=2.7u L=40.00n
.ENDS BUFV10RO_12TH40
.SUBCKT BUFV10RQ_12TH40 I Z VDD VSS
XX2 net11 I VSS VPW NHVT11LL_CKT W=680.00n L=40.00n
XX0 Z net11 VSS VPW NHVT11LL_CKT W=2.7u L=40.00n
XX1 net11 I VDD VNW PHVT11LL_CKT W=760.00n L=40.00n
XX3 Z net11 VDD VNW PHVT11LL_CKT W=3.05u L=40.00n
.ENDS BUFV10RQ_12TH40
.SUBCKT BUFV10_12TH40 I Z VDD VSS
XX2 net11 I VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX0 Z net11 VSS VPW NHVT11LL_CKT W=2.7u L=40.00n
XX1 net11 I VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX3 Z net11 VDD VNW PHVT11LL_CKT W=3.05u L=40.00n
.ENDS BUFV10_12TH40
.SUBCKT BUFV12RD_12TH40 I Z VDD VSS
XX1 net11 I VSS VPW NHVT11LL_CKT W=1.86u L=40.00n
XX6 Z net11 VSS VPW NHVT11LL_CKT W=3.24u L=40.00n
XX0 net11 I VDD VNW PHVT11LL_CKT W=2.12u L=40.00n
XX5 Z net11 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
.ENDS BUFV12RD_12TH40
.SUBCKT BUFV12RO_12TH40 I Z VDD VSS
XX1 net26 I VDD VNW PHVT11LL_CKT W=460.00n L=40.00n
XX3 Z net26 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX2 net26 I VSS VPW NHVT11LL_CKT W=405.00n L=40.00n
XX0 Z net26 VSS VPW NHVT11LL_CKT W=3.24u L=40.00n
.ENDS BUFV12RO_12TH40
.SUBCKT BUFV12RQ_12TH40 I Z VDD VSS
XX2 net11 I VSS VPW NHVT11LL_CKT W=810.00n L=40.00n
XX0 Z net11 VSS VPW NHVT11LL_CKT W=3.24u L=40.00n
XX1 net11 I VDD VNW PHVT11LL_CKT W=920.00n L=40.00n
XX3 Z net11 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
.ENDS BUFV12RQ_12TH40
.SUBCKT BUFV12_12TH40 I Z VDD VSS
XX2 net11 I VSS VPW NHVT11LL_CKT W=1.29u L=40.00n
XX0 Z net11 VSS VPW NHVT11LL_CKT W=3.21u L=40.00n
XX1 net11 I VDD VNW PHVT11LL_CKT W=1.47u L=40.00n
XX3 Z net11 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
.ENDS BUFV12_12TH40
.SUBCKT BUFV16RD_12TH40 I Z VDD VSS
XX1 net11 I VSS VPW NHVT11LL_CKT W=2.88u L=40.00n
XX6 Z net11 VSS VPW NHVT11LL_CKT W=4.32u L=40.00n
XX0 net11 I VDD VNW PHVT11LL_CKT W=3.24u L=40.00n
XX5 Z net11 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
.ENDS BUFV16RD_12TH40
.SUBCKT BUFV16RO_12TH40 I Z VDD VSS
XX1 net26 I VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX3 Z net26 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX2 net26 I VSS VPW NHVT11LL_CKT W=540.0n L=40.00n
XX0 Z net26 VSS VPW NHVT11LL_CKT W=4.32u L=40.00n
.ENDS BUFV16RO_12TH40
.SUBCKT BUFV16RQ_12TH40 I Z VDD VSS
XX2 net11 I VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX0 Z net11 VSS VPW NHVT11LL_CKT W=4.32u L=40.00n
XX1 net11 I VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX3 Z net11 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
.ENDS BUFV16RQ_12TH40
.SUBCKT BUFV16_12TH40 I Z VDD VSS
XX2 net11 I VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX0 Z net11 VSS VPW NHVT11LL_CKT W=4.32u L=40.00n
XX1 net11 I VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX3 Z net11 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
.ENDS BUFV16_12TH40
.SUBCKT BUFV1RD_12TH40 I Z VDD VSS
XX1 net11 I VSS VPW NHVT11LL_CKT W=0.265u L=40.00n
XX6 Z net11 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX0 net11 I VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX5 Z net11 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
.ENDS BUFV1RD_12TH40
.SUBCKT BUFV1_12TH40 I Z VDD VSS
XX2 net11 I VSS VPW NHVT11LL_CKT W=150.00n L=40.00n
XX0 Z net11 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX1 net11 I VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX3 Z net11 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
.ENDS BUFV1_12TH40
.SUBCKT BUFV20RD_12TH40 I Z VDD VSS
XX1 net11 I VSS VPW NHVT11LL_CKT W=3.605u L=40.00n
XX6 Z net11 VSS VPW NHVT11LL_CKT W=5.4u L=40.00n
XX0 net11 I VDD VNW PHVT11LL_CKT W=4.06u L=40.00n
XX5 Z net11 VDD VNW PHVT11LL_CKT W=6.1u L=40.00n
.ENDS BUFV20RD_12TH40
.SUBCKT BUFV20RO_12TH40 I Z VDD VSS
XX1 net26 I VDD VNW PHVT11LL_CKT W=760.00n L=40.00n
XX3 Z net26 VDD VNW PHVT11LL_CKT W=6.1u L=40.00n
XX2 net26 I VSS VPW NHVT11LL_CKT W=670.00n L=40.00n
XX0 Z net26 VSS VPW NHVT11LL_CKT W=5.4u L=40.00n
.ENDS BUFV20RO_12TH40
.SUBCKT BUFV20RQ_12TH40 I Z VDD VSS
XX2 net11 I VSS VPW NHVT11LL_CKT W=1.35u L=40.00n
XX0 Z net11 VSS VPW NHVT11LL_CKT W=5.4u L=40.00n
XX1 net11 I VDD VNW PHVT11LL_CKT W=1.53u L=40.00n
XX3 Z net11 VDD VNW PHVT11LL_CKT W=6.1u L=40.00n
.ENDS BUFV20RQ_12TH40
.SUBCKT BUFV20_12TH40 I Z VDD VSS
XX2 net11 I VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX0 Z net11 VSS VPW NHVT11LL_CKT W=5.4u L=40.00n
XX1 net11 I VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX3 Z net11 VDD VNW PHVT11LL_CKT W=6.1u L=40.00n
.ENDS BUFV20_12TH40
.SUBCKT BUFV24RD_12TH40 I Z VDD VSS
XX1 net11 I VSS VPW NHVT11LL_CKT W=4.32u L=40.00n
XX6 Z net11 VSS VPW NHVT11LL_CKT W=7.02u L=40.00n
XX0 net11 I VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX5 Z net11 VDD VNW PHVT11LL_CKT W=7.93u L=40.00n
.ENDS BUFV24RD_12TH40
.SUBCKT BUFV24RO_12TH40 I Z VDD VSS
XX1 net26 I VDD VNW PHVT11LL_CKT W=920.00n L=40.00n
XX3 Z net26 VDD VNW PHVT11LL_CKT W=7.32u L=40.00n
XX2 net26 I VSS VPW NHVT11LL_CKT W=810.00n L=40.00n
XX0 Z net26 VSS VPW NHVT11LL_CKT W=6.48u L=40.00n
.ENDS BUFV24RO_12TH40
.SUBCKT BUFV24RQ_12TH40 I Z VDD VSS
XX2 net11 I VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX0 Z net11 VSS VPW NHVT11LL_CKT W=7.02u L=40.00n
XX1 net11 I VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX3 Z net11 VDD VNW PHVT11LL_CKT W=7.93u L=40.00n
.ENDS BUFV24RQ_12TH40
.SUBCKT BUFV24_12TH40 I Z VDD VSS
XX2 net11 I VSS VPW NHVT11LL_CKT W=2.6u L=40.00n
XX0 Z net11 VSS VPW NHVT11LL_CKT W=6.48u L=40.00n
XX1 net11 I VDD VNW PHVT11LL_CKT W=2.925u L=40.00n
XX3 Z net11 VDD VNW PHVT11LL_CKT W=7.32u L=40.00n
.ENDS BUFV24_12TH40
.SUBCKT BUFV2RD_12TH40 I Z VDD VSS
XX1 net11 I VSS VPW NHVT11LL_CKT W=345.00n L=40.00n
XX6 Z net11 VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX0 net11 I VDD VNW PHVT11LL_CKT W=395.00n L=40.00n
XX5 Z net11 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS BUFV2RD_12TH40
.SUBCKT BUFV2RQ_12TH40 I Z VDD VSS
XX2 net11 I VSS VPW NHVT11LL_CKT W=135.00n L=40.00n
XX0 Z net11 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX1 net11 I VDD VNW PHVT11LL_CKT W=150.00n L=40.00n
XX3 Z net11 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS BUFV2RQ_12TH40
.SUBCKT BUFV2_12TH40 I Z VDD VSS
XX2 net11 I VSS VPW NHVT11LL_CKT W=215.00n L=40.00n
XX0 Z net11 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX1 net11 I VDD VNW PHVT11LL_CKT W=245.00n L=40.00n
XX3 Z net11 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS BUFV2_12TH40
.SUBCKT BUFV32RD_12TH40 I Z VDD VSS
XX1 net11 I VSS VPW NHVT11LL_CKT W=4.8u L=40.00n
XX6 Z net11 VSS VPW NHVT11LL_CKT W=8.64u L=40.00n
XX0 net11 I VDD VNW PHVT11LL_CKT W=5.5u L=40.00n
XX5 Z net11 VDD VNW PHVT11LL_CKT W=9.76u L=40.00n
.ENDS BUFV32RD_12TH40
.SUBCKT BUFV32RO_12TH40 I Z VDD VSS
XX1 net26 I VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX3 Z net26 VDD VNW PHVT11LL_CKT W=9.76u L=40.00n
XX2 net26 I VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX0 Z net26 VSS VPW NHVT11LL_CKT W=8.64u L=40.00n
.ENDS BUFV32RO_12TH40
.SUBCKT BUFV32RQ_12TH40 I Z VDD VSS
XX2 net11 I VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX0 Z net11 VSS VPW NHVT11LL_CKT W=8.64u L=40.00n
XX1 net11 I VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX3 Z net11 VDD VNW PHVT11LL_CKT W=9.76u L=40.00n
.ENDS BUFV32RQ_12TH40
.SUBCKT BUFV32_12TH40 I Z VDD VSS
XX2 net11 I VSS VPW NHVT11LL_CKT W=3.465u L=40.00n
XX0 Z net11 VSS VPW NHVT11LL_CKT W=8.64u L=40.00n
XX1 net11 I VDD VNW PHVT11LL_CKT W=3.92u L=40.00n
XX3 Z net11 VDD VNW PHVT11LL_CKT W=9.76u L=40.00n
.ENDS BUFV32_12TH40
.SUBCKT BUFV3RD_12TH40 I Z VDD VSS
XX1 net11 I VSS VPW NHVT11LL_CKT W=0.465u L=40.00n
XX6 Z net11 VSS VPW NHVT11LL_CKT W=0.76u L=40.00n
XX0 net11 I VDD VNW PHVT11LL_CKT W=0.53u L=40.00n
XX5 Z net11 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
.ENDS BUFV3RD_12TH40
.SUBCKT BUFV3RQ_12TH40 I Z VDD VSS
XX2 net11 I VSS VPW NHVT11LL_CKT W=190.00n L=40.00n
XX0 Z net11 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX1 net11 I VDD VNW PHVT11LL_CKT W=220.00n L=40.00n
XX3 Z net11 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
.ENDS BUFV3RQ_12TH40
.SUBCKT BUFV3_12TH40 I Z VDD VSS
XX2 net11 I VSS VPW NHVT11LL_CKT W=305.00n L=40.00n
XX0 Z net11 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX1 net11 I VDD VNW PHVT11LL_CKT W=345.00n L=40.00n
XX3 Z net11 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
.ENDS BUFV3_12TH40
.SUBCKT BUFV4RD_12TH40 I Z VDD VSS
XX1 net11 I VSS VPW NHVT11LL_CKT W=0.64u L=40.00n
XX6 Z net11 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX0 net11 I VDD VNW PHVT11LL_CKT W=0.74u L=40.00n
XX5 Z net11 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS BUFV4RD_12TH40
.SUBCKT BUFV4RO_12TH40 I Z VDD VSS
XX2 net11 I VSS VPW NHVT11LL_CKT W=135.00n L=40.00n
XX0 Z net11 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX1 net11 I VDD VNW PHVT11LL_CKT W=150.00n L=40.00n
XX3 Z net11 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS BUFV4RO_12TH40
.SUBCKT BUFV4RQ_12TH40 I Z VDD VSS
XX2 net11 I VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX0 Z net11 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX1 net11 I VDD VNW PHVT11LL_CKT W=305.00n L=40.00n
XX3 Z net11 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS BUFV4RQ_12TH40
.SUBCKT BUFV4_12TH40 I Z VDD VSS
XX2 net11 I VSS VPW NHVT11LL_CKT W=430.00n L=40.00n
XX0 Z net11 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX1 net11 I VDD VNW PHVT11LL_CKT W=490.00n L=40.00n
XX3 Z net11 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS BUFV4_12TH40
.SUBCKT BUFV5RD_12TH40 I Z VDD VSS
XX1 net11 I VSS VPW NHVT11LL_CKT W=0.79u L=40.00n
XX6 Z net11 VSS VPW NHVT11LL_CKT W=1.35u L=40.00n
XX0 net11 I VDD VNW PHVT11LL_CKT W=0.9u L=40.00n
XX5 Z net11 VDD VNW PHVT11LL_CKT W=1.53u L=40.00n
.ENDS BUFV5RD_12TH40
.SUBCKT BUFV5RO_12TH40 I Z VDD VSS
XX1 net26 I VDD VNW PHVT11LL_CKT W=190.00n L=40.00n
XX3 Z net26 VDD VNW PHVT11LL_CKT W=1.53u L=40.00n
XX2 net26 I VSS VPW NHVT11LL_CKT W=170.00n L=40.00n
XX0 Z net26 VSS VPW NHVT11LL_CKT W=1.35u L=40.00n
.ENDS BUFV5RO_12TH40
.SUBCKT BUFV5RQ_12TH40 I Z VDD VSS
XX2 net11 I VSS VPW NHVT11LL_CKT W=340.00n L=40.00n
XX0 Z net11 VSS VPW NHVT11LL_CKT W=1.35u L=40.00n
XX1 net11 I VDD VNW PHVT11LL_CKT W=380.00n L=40.00n
XX3 Z net11 VDD VNW PHVT11LL_CKT W=1.53u L=40.00n
.ENDS BUFV5RQ_12TH40
.SUBCKT BUFV5_12TH40 I Z VDD VSS
XX2 net11 I VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX0 Z net11 VSS VPW NHVT11LL_CKT W=1.35u L=40.00n
XX1 net11 I VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX3 Z net11 VDD VNW PHVT11LL_CKT W=1.53u L=40.00n
.ENDS BUFV5_12TH40
.SUBCKT BUFV6RD_12TH40 I Z VDD VSS
XX1 net11 I VSS VPW NHVT11LL_CKT W=0.92u L=40.00n
XX6 Z net11 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX0 net11 I VDD VNW PHVT11LL_CKT W=1.05u L=40.00n
XX5 Z net11 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS BUFV6RD_12TH40
.SUBCKT BUFV6RO_12TH40 I Z VDD VSS
XX1 net26 I VDD VNW PHVT11LL_CKT W=230.00n L=40.00n
XX3 Z net26 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX2 net26 I VSS VPW NHVT11LL_CKT W=200.00n L=40.00n
XX0 Z net26 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
.ENDS BUFV6RO_12TH40
.SUBCKT BUFV6RQ_12TH40 I Z VDD VSS
XX2 net11 I VSS VPW NHVT11LL_CKT W=405.00n L=40.00n
XX0 Z net11 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX1 net11 I VDD VNW PHVT11LL_CKT W=460.00n L=40.00n
XX3 Z net11 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS BUFV6RQ_12TH40
.SUBCKT BUFV6_12TH40 I Z VDD VSS
XX2 net11 I VSS VPW NHVT11LL_CKT W=650.00n L=40.00n
XX0 Z net11 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX1 net11 I VDD VNW PHVT11LL_CKT W=730.00n L=40.00n
XX3 Z net11 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS BUFV6_12TH40
.SUBCKT BUFV7RD_12TH40 I Z VDD VSS
XX1 net11 I VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX6 Z net11 VSS VPW NHVT11LL_CKT W=1.88u L=40.00n
XX0 net11 I VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX5 Z net11 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
.ENDS BUFV7RD_12TH40
.SUBCKT BUFV7RO_12TH40 I Z VDD VSS
XX1 net26 I VDD VNW PHVT11LL_CKT W=270.00n L=40.00n
XX3 Z net26 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
XX2 net26 I VSS VPW NHVT11LL_CKT W=235.00n L=40.00n
XX0 Z net26 VSS VPW NHVT11LL_CKT W=1.88u L=40.00n
.ENDS BUFV7RO_12TH40
.SUBCKT BUFV7RQ_12TH40 I Z VDD VSS
XX2 net11 I VSS VPW NHVT11LL_CKT W=470.00n L=40.00n
XX0 Z net11 VSS VPW NHVT11LL_CKT W=1.88u L=40.00n
XX1 net11 I VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX3 Z net11 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
.ENDS BUFV7RQ_12TH40
.SUBCKT BUFV7_12TH40 I Z VDD VSS
XX2 net11 I VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX0 Z net11 VSS VPW NHVT11LL_CKT W=1.88u L=40.00n
XX1 net11 I VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX3 Z net11 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
.ENDS BUFV7_12TH40
.SUBCKT BUFV8RD_12TH40 I Z VDD VSS
XX1 net11 I VSS VPW NHVT11LL_CKT W=1.26u L=40.00n
XX6 Z net11 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX0 net11 I VDD VNW PHVT11LL_CKT W=1.44u L=40.00n
XX5 Z net11 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS BUFV8RD_12TH40
.SUBCKT BUFV8RO_12TH40 I Z VDD VSS
XX1 net26 I VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
XX3 Z net26 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX2 net26 I VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX0 Z net26 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
.ENDS BUFV8RO_12TH40
.SUBCKT BUFV8RQ_12TH40 I Z VDD VSS
XX2 net11 I VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX0 Z net11 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX1 net11 I VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX3 Z net11 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS BUFV8RQ_12TH40
.SUBCKT BUFV8_12TH40 I Z VDD VSS
XX2 net11 I VSS VPW NHVT11LL_CKT W=860.00n L=40.00n
XX0 Z net11 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX1 net11 I VDD VNW PHVT11LL_CKT W=980.00n L=40.00n
XX3 Z net11 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS BUFV8_12TH40
.SUBCKT CLKAND2V0_12TH40 A1 A2 Z VDD VSS
XX6 Z net026 VSS VPW NHVT11LL_CKT W=130.00n L=40.00n
XX9 net026 A1 net4 VPW NHVT11LL_CKT W=130.00n L=40.00n
XX8 net4 A2 VSS VPW NHVT11LL_CKT W=130.00n L=40.00n
XX5 Z net026 VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
XX28 net026 A1 VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX0 net026 A2 VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
.ENDS CLKAND2V0_12TH40
.SUBCKT CLKAND2V12_12TH40 A1 A2 Z VDD VSS
XX6 Z net026 VSS VPW NHVT11LL_CKT W=1.56u L=40.00n
XX9 net026 A1 net4 VPW NHVT11LL_CKT W=960.00n L=40.00n
XX8 net4 A2 VSS VPW NHVT11LL_CKT W=960.00n L=40.00n
XX5 Z net026 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX28 net026 A1 VDD VNW PHVT11LL_CKT W=1.03u L=40.00n
XX0 net026 A2 VDD VNW PHVT11LL_CKT W=1.03u L=40.00n
.ENDS CLKAND2V12_12TH40
.SUBCKT CLKAND2V16_12TH40 A1 A2 Z VDD VSS
XX6 Z net026 VSS VPW NHVT11LL_CKT W=2.08u L=40.00n
XX9 net026 A1 net4 VPW NHVT11LL_CKT W=1.35u L=40.00n
XX8 net4 A2 VSS VPW NHVT11LL_CKT W=1.35u L=40.00n
XX5 Z net026 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX28 net026 A1 VDD VNW PHVT11LL_CKT W=1.47u L=40.00n
XX0 net026 A2 VDD VNW PHVT11LL_CKT W=1.47u L=40.00n
.ENDS CLKAND2V16_12TH40
.SUBCKT CLKAND2V1_12TH40 A1 A2 Z VDD VSS
XX6 Z net026 VSS VPW NHVT11LL_CKT W=185.00n L=40.00n
XX9 net026 A1 net4 VPW NHVT11LL_CKT W=165.00n L=40.00n
XX8 net4 A2 VSS VPW NHVT11LL_CKT W=165.00n L=40.00n
XX5 Z net026 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX28 net026 A1 VDD VNW PHVT11LL_CKT W=185.00n L=40.00n
XX0 net026 A2 VDD VNW PHVT11LL_CKT W=185.00n L=40.00n
.ENDS CLKAND2V1_12TH40
.SUBCKT CLKAND2V20_12TH40 A1 A2 Z VDD VSS
XX6 Z net026 VSS VPW NHVT11LL_CKT W=2.6u L=40.00n
XX9 net026 A1 net4 VPW NHVT11LL_CKT W=1.665u L=40.00n
XX8 net4 A2 VSS VPW NHVT11LL_CKT W=1.665u L=40.00n
XX5 Z net026 VDD VNW PHVT11LL_CKT W=6.1u L=40.00n
XX28 net026 A1 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX0 net026 A2 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS CLKAND2V20_12TH40
.SUBCKT CLKAND2V24_12TH40 A1 A2 Z VDD VSS
XX6 Z net026 VSS VPW NHVT11LL_CKT W=3.12u L=40.00n
XX9 net026 A1 net4 VPW NHVT11LL_CKT W=2.22u L=40.00n
XX8 net4 A2 VSS VPW NHVT11LL_CKT W=2.22u L=40.00n
XX5 Z net026 VDD VNW PHVT11LL_CKT W=7.32u L=40.00n
XX28 net026 A1 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX0 net026 A2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS CLKAND2V24_12TH40
.SUBCKT CLKAND2V2_12TH40 A1 A2 Z VDD VSS
XX6 Z net026 VSS VPW NHVT11LL_CKT W=260.00n L=40.00n
XX9 net026 A1 net4 VPW NHVT11LL_CKT W=190.00n L=40.00n
XX8 net4 A2 VSS VPW NHVT11LL_CKT W=190.00n L=40.00n
XX5 Z net026 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX28 net026 A1 VDD VNW PHVT11LL_CKT W=210.00n L=40.00n
XX0 net026 A2 VDD VNW PHVT11LL_CKT W=210.00n L=40.00n
.ENDS CLKAND2V2_12TH40
.SUBCKT CLKAND2V3_12TH40 A1 A2 Z VDD VSS
XX6 Z net026 VSS VPW NHVT11LL_CKT W=370.00n L=40.00n
XX9 net026 A1 net4 VPW NHVT11LL_CKT W=255.00n L=40.00n
XX8 net4 A2 VSS VPW NHVT11LL_CKT W=255.00n L=40.00n
XX5 Z net026 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX28 net026 A1 VDD VNW PHVT11LL_CKT W=280.00n L=40.00n
XX0 net026 A2 VDD VNW PHVT11LL_CKT W=280.00n L=40.00n
.ENDS CLKAND2V3_12TH40
.SUBCKT CLKAND2V4_12TH40 A1 A2 Z VDD VSS
XX6 Z net026 VSS VPW NHVT11LL_CKT W=520.00n L=40.00n
XX9 net026 A1 net4 VPW NHVT11LL_CKT W=345.00n L=40.00n
XX8 net4 A2 VSS VPW NHVT11LL_CKT W=345.00n L=40.00n
XX5 Z net026 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX28 net026 A1 VDD VNW PHVT11LL_CKT W=380.00n L=40.00n
XX0 net026 A2 VDD VNW PHVT11LL_CKT W=380.00n L=40.00n
.ENDS CLKAND2V4_12TH40
.SUBCKT CLKAND2V6_12TH40 A1 A2 Z VDD VSS
XX6 Z net026 VSS VPW NHVT11LL_CKT W=780.00n L=40.00n
XX9 net026 A1 net4 VPW NHVT11LL_CKT W=480.00n L=40.00n
XX8 net4 A2 VSS VPW NHVT11LL_CKT W=480.00n L=40.00n
XX5 Z net026 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX28 net026 A1 VDD VNW PHVT11LL_CKT W=530.00n L=40.00n
XX0 net026 A2 VDD VNW PHVT11LL_CKT W=530.00n L=40.00n
.ENDS CLKAND2V6_12TH40
.SUBCKT CLKAND2V8_12TH40 A1 A2 Z VDD VSS
XX6 Z net026 VSS VPW NHVT11LL_CKT W=1.04u L=40.00n
XX9 net026 A1 net4 VPW NHVT11LL_CKT W=670.00n L=40.00n
XX8 net4 A2 VSS VPW NHVT11LL_CKT W=670.00n L=40.00n
XX5 Z net026 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX28 net026 A1 VDD VNW PHVT11LL_CKT W=740.00n L=40.00n
XX0 net026 A2 VDD VNW PHVT11LL_CKT W=740.00n L=40.00n
.ENDS CLKAND2V8_12TH40
.SUBCKT CLKBUFV10RQ_12TH40 I Z VDD VSS
XX0 Z net7 VSS VPW NHVT11LL_CKT W=1.3u L=40.00n
XX2 net7 I VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX3 Z net7 VDD VNW PHVT11LL_CKT W=3.05u L=40.00n
XX1 net7 I VDD VNW PHVT11LL_CKT W=760.00n L=40.00n
.ENDS CLKBUFV10RQ_12TH40
.SUBCKT CLKBUFV10_12TH40 I Z VDD VSS
XX0 Z net7 VSS VPW NHVT11LL_CKT W=1.3u L=40.00n
XX2 net7 I VSS VPW NHVT11LL_CKT W=520.00n L=40.00n
XX3 Z net7 VDD VNW PHVT11LL_CKT W=3.05u L=40.00n
XX1 net7 I VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS CLKBUFV10_12TH40
.SUBCKT CLKBUFV12RQ_12TH40 I Z VDD VSS
XX0 Z net7 VSS VPW NHVT11LL_CKT W=1.56u L=40.00n
XX2 net7 I VSS VPW NHVT11LL_CKT W=390.00n L=40.00n
XX3 Z net7 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX1 net7 I VDD VNW PHVT11LL_CKT W=920.00n L=40.00n
.ENDS CLKBUFV12RQ_12TH40
.SUBCKT CLKBUFV12_12TH40 I Z VDD VSS
XX0 Z net7 VSS VPW NHVT11LL_CKT W=1.56u L=40.00n
XX2 net7 I VSS VPW NHVT11LL_CKT W=630.00n L=40.00n
XX3 Z net7 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX1 net7 I VDD VNW PHVT11LL_CKT W=1.47u L=40.00n
.ENDS CLKBUFV12_12TH40
.SUBCKT CLKBUFV16RQ_12TH40 I Z VDD VSS
XX0 Z net7 VSS VPW NHVT11LL_CKT W=2.08u L=40.00n
XX2 net7 I VSS VPW NHVT11LL_CKT W=520.00n L=40.00n
XX3 Z net7 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX1 net7 I VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS CLKBUFV16RQ_12TH40
.SUBCKT CLKBUFV16_12TH40 I Z VDD VSS
XX0 Z net7 VSS VPW NHVT11LL_CKT W=2.08u L=40.00n
XX2 net7 I VSS VPW NHVT11LL_CKT W=780.00n L=40.00n
XX3 Z net7 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX1 net7 I VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS CLKBUFV16_12TH40
.SUBCKT CLKBUFV1_12TH40 I Z VDD VSS
XX0 Z net7 VSS VPW NHVT11LL_CKT W=185.00n L=40.00n
XX2 net7 I VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX3 Z net7 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX1 net7 I VDD VNW PHVT11LL_CKT W=280.00n L=40.00n
.ENDS CLKBUFV1_12TH40
.SUBCKT CLKBUFV20RQ_12TH40 I Z VDD VSS
XX0 Z net7 VSS VPW NHVT11LL_CKT W=2.6u L=40.00n
XX2 net7 I VSS VPW NHVT11LL_CKT W=660.00n L=40.00n
XX3 Z net7 VDD VNW PHVT11LL_CKT W=6.1u L=40.00n
XX1 net7 I VDD VNW PHVT11LL_CKT W=1.53u L=40.00n
.ENDS CLKBUFV20RQ_12TH40
.SUBCKT CLKBUFV20_12TH40 I Z VDD VSS
XX0 Z net7 VSS VPW NHVT11LL_CKT W=2.6u L=40.00n
XX2 net7 I VSS VPW NHVT11LL_CKT W=1.04u L=40.00n
XX3 Z net7 VDD VNW PHVT11LL_CKT W=6.1u L=40.00n
XX1 net7 I VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS CLKBUFV20_12TH40
.SUBCKT CLKBUFV24RQ_12TH40 I Z VDD VSS
XX0 Z net7 VSS VPW NHVT11LL_CKT W=3.12u L=40.00n
XX2 net7 I VSS VPW NHVT11LL_CKT W=780.00n L=40.00n
XX3 Z net7 VDD VNW PHVT11LL_CKT W=7.32u L=40.00n
XX1 net7 I VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS CLKBUFV24RQ_12TH40
.SUBCKT CLKBUFV24_12TH40 I Z VDD VSS
XX0 Z net7 VSS VPW NHVT11LL_CKT W=3.12u L=40.00n
XX2 net7 I VSS VPW NHVT11LL_CKT W=1.3u L=40.00n
XX3 Z net7 VDD VNW PHVT11LL_CKT W=7.32u L=40.00n
XX1 net7 I VDD VNW PHVT11LL_CKT W=3.05u L=40.00n
.ENDS CLKBUFV24_12TH40
.SUBCKT CLKBUFV2_12TH40 I Z VDD VSS
XX0 Z net7 VSS VPW NHVT11LL_CKT W=260.00n L=40.00n
XX2 net7 I VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX3 Z net7 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 net7 I VDD VNW PHVT11LL_CKT W=280.00n L=40.00n
.ENDS CLKBUFV2_12TH40
.SUBCKT CLKBUFV32_12TH40 I Z VDD VSS
XX0 Z net7 VSS VPW NHVT11LL_CKT W=4.16u L=40.00n
XX2 net7 I VSS VPW NHVT11LL_CKT W=1.68u L=40.00n
XX3 Z net7 VDD VNW PHVT11LL_CKT W=9.76u L=40.00n
XX1 net7 I VDD VNW PHVT11LL_CKT W=3.92u L=40.00n
.ENDS CLKBUFV32_12TH40
.SUBCKT CLKBUFV3_12TH40 I Z VDD VSS
XX0 Z net7 VSS VPW NHVT11LL_CKT W=370.00n L=40.00n
XX2 net7 I VSS VPW NHVT11LL_CKT W=145.00n L=40.00n
XX3 Z net7 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX1 net7 I VDD VNW PHVT11LL_CKT W=345.00n L=40.00n
.ENDS CLKBUFV3_12TH40
.SUBCKT CLKBUFV4RQ_12TH40 I Z VDD VSS
XX0 Z net7 VSS VPW NHVT11LL_CKT W=520.00n L=40.00n
XX2 net7 I VSS VPW NHVT11LL_CKT W=130.00n L=40.00n
XX3 Z net7 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 net7 I VDD VNW PHVT11LL_CKT W=305.00n L=40.00n
.ENDS CLKBUFV4RQ_12TH40
.SUBCKT CLKBUFV4_12TH40 I Z VDD VSS
XX0 Z net7 VSS VPW NHVT11LL_CKT W=520.00n L=40.00n
XX2 net7 I VSS VPW NHVT11LL_CKT W=210.00n L=40.00n
XX3 Z net7 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 net7 I VDD VNW PHVT11LL_CKT W=490.00n L=40.00n
.ENDS CLKBUFV4_12TH40
.SUBCKT CLKBUFV5_12TH40 I Z VDD VSS
XX0 Z net7 VSS VPW NHVT11LL_CKT W=650.00n L=40.00n
XX2 net7 I VSS VPW NHVT11LL_CKT W=260.00n L=40.00n
XX3 Z net7 VDD VNW PHVT11LL_CKT W=1.53u L=40.00n
XX1 net7 I VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS CLKBUFV5_12TH40
.SUBCKT CLKBUFV6RQ_12TH40 I Z VDD VSS
XX0 Z net7 VSS VPW NHVT11LL_CKT W=780.00n L=40.00n
XX2 net7 I VSS VPW NHVT11LL_CKT W=195.00n L=40.00n
XX3 Z net7 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX1 net7 I VDD VNW PHVT11LL_CKT W=460.00n L=40.00n
.ENDS CLKBUFV6RQ_12TH40
.SUBCKT CLKBUFV6_12TH40 I Z VDD VSS
XX0 Z net7 VSS VPW NHVT11LL_CKT W=780.00n L=40.00n
XX2 net7 I VSS VPW NHVT11LL_CKT W=310.00n L=40.00n
XX3 Z net7 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX1 net7 I VDD VNW PHVT11LL_CKT W=730.00n L=40.00n
.ENDS CLKBUFV6_12TH40
.SUBCKT CLKBUFV7_12TH40 I Z VDD VSS
XX0 Z net7 VSS VPW NHVT11LL_CKT W=920.00n L=40.00n
XX2 net7 I VSS VPW NHVT11LL_CKT W=370.00n L=40.00n
XX3 Z net7 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
XX1 net7 I VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
.ENDS CLKBUFV7_12TH40
.SUBCKT CLKBUFV8RQ_12TH40 I Z VDD VSS
XX0 Z net7 VSS VPW NHVT11LL_CKT W=1.04u L=40.00n
XX2 net7 I VSS VPW NHVT11LL_CKT W=260.00n L=40.00n
XX3 Z net7 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 net7 I VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS CLKBUFV8RQ_12TH40
.SUBCKT CLKBUFV8_12TH40 I Z VDD VSS
XX0 Z net7 VSS VPW NHVT11LL_CKT W=1.04u L=40.00n
XX2 net7 I VSS VPW NHVT11LL_CKT W=420.00n L=40.00n
XX3 Z net7 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 net7 I VDD VNW PHVT11LL_CKT W=980.00n L=40.00n
.ENDS CLKBUFV8_12TH40
.SUBCKT CLKINV0_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=130.00n L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
.ENDS CLKINV0_12TH40
.SUBCKT CLKINV10_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=1.3u L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=3.05u L=40.00n
.ENDS CLKINV10_12TH40
.SUBCKT CLKINV12_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=1.56u L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
.ENDS CLKINV12_12TH40
.SUBCKT CLKINV16_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=2.08u L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
.ENDS CLKINV16_12TH40
.SUBCKT CLKINV1_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=185.00n L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
.ENDS CLKINV1_12TH40
.SUBCKT CLKINV20_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=2.6u L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=6.1u L=40.00n
.ENDS CLKINV20_12TH40
.SUBCKT CLKINV24_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=3.12u L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=7.32u L=40.00n
.ENDS CLKINV24_12TH40
.SUBCKT CLKINV2_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=260.00n L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS CLKINV2_12TH40
.SUBCKT CLKINV32_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=4.16u L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=9.76u L=40.00n
.ENDS CLKINV32_12TH40
.SUBCKT CLKINV3_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=370.00n L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
.ENDS CLKINV3_12TH40
.SUBCKT CLKINV4_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=520.00n L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS CLKINV4_12TH40
.SUBCKT CLKINV5_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=650.00n L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=1.53u L=40.00n
.ENDS CLKINV5_12TH40
.SUBCKT CLKINV6_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=780.00n L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS CLKINV6_12TH40
.SUBCKT CLKINV7_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=920.00n L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
.ENDS CLKINV7_12TH40
.SUBCKT CLKINV8_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=1.04u L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS CLKINV8_12TH40
.SUBCKT CLKLAHAQV0_12TH40 CK E Q TE VDD VSS
XX20 ten TE VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX15 Q s VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
XX16 nt11 E VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX17 pm cn nt11 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX18 cn CK VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX13 nt21 pm VDD VNW PHVT11LL_CKT W=560.00n L=40.00n
XX14 s CK nt21 VNW PHVT11LL_CKT W=560.00n L=40.00n
XX21 m pm VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX12 nt21 ten VDD VNW PHVT11LL_CKT W=560.00n L=40.00n
XX22 nt13 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 pm CK nt13 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 ten TE VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX1 nt12 E VSS VPW NHVT11LL_CKT W=0.24u L=40.00n
XX3 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX9 nt22 ten VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX10 pm cn nt14 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 Q s VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX6 s pm nt22 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX0 pm CK nt12 VPW NHVT11LL_CKT W=0.24u L=40.00n
XX2 m pm VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX8 s CK VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX11 nt14 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
.ENDS CLKLAHAQV0_12TH40
.SUBCKT CLKLAHAQV10_12TH40 CK E Q TE VDD VSS
XX20 ten TE VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX15 Q s VDD VNW PHVT11LL_CKT W=3.05u L=40.00n
XX16 nt11 E VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX17 pm cn nt11 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX18 cn CK VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX13 nt21 pm VDD VNW PHVT11LL_CKT W=1.04u L=40.00n
XX14 s CK nt21 VNW PHVT11LL_CKT W=1.04u L=40.00n
XX21 m pm VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX12 nt21 ten VDD VNW PHVT11LL_CKT W=1.04u L=40.00n
XX22 nt13 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 pm CK nt13 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 ten TE VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX1 nt12 E VSS VPW NHVT11LL_CKT W=0.335u L=40.00n
XX3 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX9 nt22 ten VSS VPW NHVT11LL_CKT W=240.00n L=40.00n
XX10 pm cn nt14 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 Q s VSS VPW NHVT11LL_CKT W=1.3u L=40.00n
XX6 s pm nt22 VPW NHVT11LL_CKT W=240.00n L=40.00n
XX0 pm CK nt12 VPW NHVT11LL_CKT W=0.335u L=40.00n
XX2 m pm VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX8 s CK VSS VPW NHVT11LL_CKT W=240.00n L=40.00n
XX11 nt14 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
.ENDS CLKLAHAQV10_12TH40
.SUBCKT CLKLAHAQV12_12TH40 CK E Q TE VDD VSS
XX20 ten TE VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX15 Q s VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX16 nt11 E VDD VNW PHVT11LL_CKT W=0.52u L=40.00n
XX17 pm cn nt11 VNW PHVT11LL_CKT W=0.52u L=40.00n
XX18 cn CK VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX13 nt21 pm VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX14 s CK nt21 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX21 m pm VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX12 nt21 ten VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX22 nt13 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 pm CK nt13 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 ten TE VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX1 nt12 E VSS VPW NHVT11LL_CKT W=0.345u L=40.00n
XX3 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX9 nt22 ten VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX10 pm cn nt14 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 Q s VSS VPW NHVT11LL_CKT W=1.56u L=40.00n
XX6 s pm nt22 VPW NHVT11LL_CKT W=0.27u L=40.00n
XX0 pm CK nt12 VPW NHVT11LL_CKT W=0.345u L=40.00n
XX2 m pm VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX8 s CK VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX11 nt14 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
.ENDS CLKLAHAQV12_12TH40
.SUBCKT CLKLAHAQV16_12TH40 CK E Q TE VDD VSS
XX20 ten TE VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX15 Q s VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX16 nt11 E VDD VNW PHVT11LL_CKT W=0.55u L=40.00n
XX17 pm cn nt11 VNW PHVT11LL_CKT W=0.55u L=40.00n
XX18 cn CK VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX13 nt21 pm VDD VNW PHVT11LL_CKT W=1.5u L=40.00n
XX14 s CK nt21 VNW PHVT11LL_CKT W=1.5u L=40.00n
XX21 m pm VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX12 nt21 ten VDD VNW PHVT11LL_CKT W=1.5u L=40.00n
XX22 nt13 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 pm CK nt13 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 ten TE VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX1 nt12 E VSS VPW NHVT11LL_CKT W=0.365u L=40.00n
XX3 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX9 nt22 ten VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX10 pm cn nt14 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 Q s VSS VPW NHVT11LL_CKT W=2.08u L=40.00n
XX6 s pm nt22 VPW NHVT11LL_CKT W=380.00n L=40.00n
XX0 pm CK nt12 VPW NHVT11LL_CKT W=0.365u L=40.00n
XX2 m pm VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX8 s CK VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX11 nt14 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
.ENDS CLKLAHAQV16_12TH40
.SUBCKT CLKLAHAQV1_12TH40 CK E Q TE VDD VSS
XX20 ten TE VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX15 Q s VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX16 nt11 E VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX17 pm cn nt11 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX18 cn CK VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX13 nt21 pm VDD VNW PHVT11LL_CKT W=0.58u L=40.00n
XX14 s CK nt21 VNW PHVT11LL_CKT W=0.58u L=40.00n
XX21 m pm VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX12 nt21 ten VDD VNW PHVT11LL_CKT W=0.58u L=40.00n
XX22 nt13 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 pm CK nt13 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 ten TE VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX1 nt12 E VSS VPW NHVT11LL_CKT W=0.24u L=40.00n
XX3 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX9 nt22 ten VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX10 pm cn nt14 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 Q s VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX6 s pm nt22 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX0 pm CK nt12 VPW NHVT11LL_CKT W=0.24u L=40.00n
XX2 m pm VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX8 s CK VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX11 nt14 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
.ENDS CLKLAHAQV1_12TH40
.SUBCKT CLKLAHAQV20_12TH40 CK E Q TE VDD VSS
XX20 ten TE VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX15 Q s VDD VNW PHVT11LL_CKT W=6.1u L=40.00n
XX16 nt11 E VDD VNW PHVT11LL_CKT W=0.58u L=40.00n
XX17 pm cn nt11 VNW PHVT11LL_CKT W=0.58u L=40.00n
XX18 cn CK VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX13 nt21 pm VDD VNW PHVT11LL_CKT W=1.65u L=40.00n
XX14 s CK nt21 VNW PHVT11LL_CKT W=1.65u L=40.00n
XX21 m pm VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX12 nt21 ten VDD VNW PHVT11LL_CKT W=1.65u L=40.00n
XX22 nt13 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 pm CK nt13 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 ten TE VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX1 nt12 E VSS VPW NHVT11LL_CKT W=0.385u L=40.00n
XX3 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX9 nt22 ten VSS VPW NHVT11LL_CKT W=0.36u L=40.00n
XX10 pm cn nt14 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 Q s VSS VPW NHVT11LL_CKT W=2.6u L=40.00n
XX6 s pm nt22 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX0 pm CK nt12 VPW NHVT11LL_CKT W=0.385u L=40.00n
XX2 m pm VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX8 s CK VSS VPW NHVT11LL_CKT W=0.36u L=40.00n
XX11 nt14 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
.ENDS CLKLAHAQV20_12TH40
.SUBCKT CLKLAHAQV24_12TH40 CK E Q TE VDD VSS
XX5 ten TE VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX1 nt12 E VSS VPW NHVT11LL_CKT W=0.405u L=40.00n
XX3 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX9 nt22 ten VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX10 pm cn nt14 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 Q s VSS VPW NHVT11LL_CKT W=3.12u L=40.00n
XX6 s pm nt22 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX0 pm CK nt12 VPW NHVT11LL_CKT W=0.405u L=40.00n
XX2 m pm VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX8 s CK VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX11 nt14 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX20 ten TE VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX15 Q s VDD VNW PHVT11LL_CKT W=7.32u L=40.00n
XX16 nt11 E VDD VNW PHVT11LL_CKT W=0.595u L=40.00n
XX17 pm cn nt11 VNW PHVT11LL_CKT W=0.595u L=40.00n
XX18 cn CK VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX13 nt21 pm VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX14 s CK nt21 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX21 m pm VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX12 nt21 ten VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX22 nt13 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 pm CK nt13 VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS CLKLAHAQV24_12TH40
.SUBCKT CLKLAHAQV2_12TH40 CK E Q TE VDD VSS
XX20 ten TE VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX15 Q s VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX16 nt11 E VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX17 pm cn nt11 VNW PHVT11LL_CKT W=0.4u L=40.00n
XX18 cn CK VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX13 nt21 pm VDD VNW PHVT11LL_CKT W=0.59u L=40.00n
XX14 s CK nt21 VNW PHVT11LL_CKT W=0.59u L=40.00n
XX21 m pm VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX12 nt21 ten VDD VNW PHVT11LL_CKT W=0.59u L=40.00n
XX22 nt13 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 pm CK nt13 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 ten TE VSS VPW NHVT11LL_CKT W=170.00n L=40.00n
XX1 nt12 E VSS VPW NHVT11LL_CKT W=0.26u L=40.00n
XX3 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX9 nt22 ten VSS VPW NHVT11LL_CKT W=140.00n L=40.00n
XX10 pm cn nt14 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 Q s VSS VPW NHVT11LL_CKT W=0.26u L=40.00n
XX6 s pm nt22 VPW NHVT11LL_CKT W=140.00n L=40.00n
XX0 pm CK nt12 VPW NHVT11LL_CKT W=0.26u L=40.00n
XX2 m pm VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX8 s CK VSS VPW NHVT11LL_CKT W=140.00n L=40.00n
XX11 nt14 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
.ENDS CLKLAHAQV2_12TH40
.SUBCKT CLKLAHAQV3_12TH40 CK E Q TE VDD VSS
XX20 ten TE VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX15 Q s VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX16 nt11 E VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX17 pm cn nt11 VNW PHVT11LL_CKT W=0.42u L=40.00n
XX18 cn CK VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX13 nt21 pm VDD VNW PHVT11LL_CKT W=0.68u L=40.00n
XX14 s CK nt21 VNW PHVT11LL_CKT W=0.68u L=40.00n
XX21 m pm VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX12 nt21 ten VDD VNW PHVT11LL_CKT W=0.68u L=40.00n
XX22 nt13 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 pm CK nt13 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 ten TE VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX1 nt12 E VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX3 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX9 nt22 ten VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX10 pm cn nt14 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 Q s VSS VPW NHVT11LL_CKT W=0.37u L=40.00n
XX6 s pm nt22 VPW NHVT11LL_CKT W=0.16u L=40.00n
XX0 pm CK nt12 VPW NHVT11LL_CKT W=0.28u L=40.00n
XX2 m pm VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX8 s CK VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX11 nt14 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
.ENDS CLKLAHAQV3_12TH40
.SUBCKT CLKLAHAQV4_12TH40 CK E Q TE VDD VSS
XX20 ten TE VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX15 Q s VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX16 nt11 E VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX17 pm cn nt11 VNW PHVT11LL_CKT W=0.44u L=40.00n
XX18 cn CK VDD VNW PHVT11LL_CKT W=0.26u L=40.00n
XX13 nt21 pm VDD VNW PHVT11LL_CKT W=0.74u L=40.00n
XX14 s CK nt21 VNW PHVT11LL_CKT W=0.74u L=40.00n
XX21 m pm VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX12 nt21 ten VDD VNW PHVT11LL_CKT W=0.74u L=40.00n
XX22 nt13 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 pm CK nt13 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 ten TE VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX1 nt12 E VSS VPW NHVT11LL_CKT W=0.295u L=40.00n
XX3 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX9 nt22 ten VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX10 pm cn nt14 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 Q s VSS VPW NHVT11LL_CKT W=0.52u L=40.00n
XX6 s pm nt22 VPW NHVT11LL_CKT W=0.16u L=40.00n
XX0 pm CK nt12 VPW NHVT11LL_CKT W=0.295u L=40.00n
XX2 m pm VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX8 s CK VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX11 nt14 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
.ENDS CLKLAHAQV4_12TH40
.SUBCKT CLKLAHAQV6_12TH40 CK E Q TE VDD VSS
XX20 ten TE VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX15 Q s VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX16 nt11 E VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
XX17 pm cn nt11 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX18 cn CK VDD VNW PHVT11LL_CKT W=0.26u L=40.00n
XX13 nt21 pm VDD VNW PHVT11LL_CKT W=0.84u L=40.00n
XX14 s CK nt21 VNW PHVT11LL_CKT W=0.84u L=40.00n
XX21 m pm VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX12 nt21 ten VDD VNW PHVT11LL_CKT W=0.84u L=40.00n
XX22 nt13 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 pm CK nt13 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 ten TE VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX1 nt12 E VSS VPW NHVT11LL_CKT W=0.305u L=40.00n
XX3 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX9 nt22 ten VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX10 pm cn nt14 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 Q s VSS VPW NHVT11LL_CKT W=0.78u L=40.00n
XX6 s pm nt22 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX0 pm CK nt12 VPW NHVT11LL_CKT W=0.305u L=40.00n
XX2 m pm VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX8 s CK VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX11 nt14 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
.ENDS CLKLAHAQV6_12TH40
.SUBCKT CLKLAHAQV8_12TH40 CK E Q TE VDD VSS
XX20 ten TE VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX15 Q s VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX16 nt11 E VDD VNW PHVT11LL_CKT W=0.48u L=40.00n
XX17 pm cn nt11 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX18 cn CK VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX13 nt21 pm VDD VNW PHVT11LL_CKT W=1.00u L=40.00n
XX14 s CK nt21 VNW PHVT11LL_CKT W=1.00u L=40.00n
XX21 m pm VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX12 nt21 ten VDD VNW PHVT11LL_CKT W=1.00u L=40.00n
XX22 nt13 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 pm CK nt13 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 ten TE VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX1 nt12 E VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX3 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX9 nt22 ten VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX10 pm cn nt14 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 Q s VSS VPW NHVT11LL_CKT W=1.04u L=40.00n
XX6 s pm nt22 VPW NHVT11LL_CKT W=0.23u L=40.00n
XX0 pm CK nt12 VPW NHVT11LL_CKT W=0.32u L=40.00n
XX2 m pm VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX8 s CK VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX11 nt14 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
.ENDS CLKLAHAQV8_12TH40
.SUBCKT CLKLAHQV0_12TH40 CK E Q TE VDD VSS
XX6 hnet31 pm VDD VNW PHVT11LL_CKT W=0.57u L=40.00n
XX7 s CK hnet31 VNW PHVT11LL_CKT W=0.57u L=40.00n
XX9 hnet21 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX2 hnet13 TE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX3 hnet11 E hnet13 VNW PHVT11LL_CKT W=0.395u L=40.00n
XX5 m pm VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX10 pm CK hnet21 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 Q s VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
XX4 pm cn hnet11 VNW PHVT11LL_CKT W=0.395u L=40.00n
XX0 cn CK VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX20 pm cn hnet22 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 hnet12 TE VSS VPW NHVT11LL_CKT W=200.00n L=40.00n
XX15 hnet12 E VSS VPW NHVT11LL_CKT W=200.00n L=40.00n
XX16 m pm VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX19 Q s VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX13 pm CK hnet12 VPW NHVT11LL_CKT W=200.00n L=40.00n
XX18 s CK VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX11 cn CK VSS VPW NHVT11LL_CKT W=170.00n L=40.00n
XX17 s pm VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX21 hnet22 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
.ENDS CLKLAHQV0_12TH40
.SUBCKT CLKLAHQV10_12TH40 CK E Q TE VDD VSS
XX6 hnet31 pm VDD VNW PHVT11LL_CKT W=1.1u L=40.00n
XX7 s CK hnet31 VNW PHVT11LL_CKT W=1.1u L=40.00n
XX9 hnet21 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX2 hnet13 TE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX3 hnet11 E hnet13 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX5 m pm VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX10 pm CK hnet21 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 Q s VDD VNW PHVT11LL_CKT W=3.05u L=40.00n
XX4 pm cn hnet11 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 cn CK VDD VNW PHVT11LL_CKT W=0.18u L=40.00n
XX20 pm cn hnet22 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 hnet12 TE VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX15 hnet12 E VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX16 m pm VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX19 Q s VSS VPW NHVT11LL_CKT W=1.3u L=40.00n
XX13 pm CK hnet12 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX18 s CK VSS VPW NHVT11LL_CKT W=0.26u L=40.00n
XX11 cn CK VSS VPW NHVT11LL_CKT W=170.00n L=40.00n
XX17 s pm VSS VPW NHVT11LL_CKT W=0.26u L=40.00n
XX21 hnet22 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
.ENDS CLKLAHQV10_12TH40
.SUBCKT CLKLAHQV12_12TH40 CK E Q TE VDD VSS
XX6 hnet31 pm VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX7 s CK hnet31 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX9 hnet21 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX2 hnet13 TE VDD VNW PHVT11LL_CKT W=0.8u L=40.00n
XX3 hnet11 E hnet13 VNW PHVT11LL_CKT W=0.8u L=40.00n
XX5 m pm VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX10 pm CK hnet21 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 Q s VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX4 pm cn hnet11 VNW PHVT11LL_CKT W=0.8u L=40.00n
XX0 cn CK VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX20 pm cn hnet22 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 hnet12 TE VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX15 hnet12 E VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX16 m pm VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX19 Q s VSS VPW NHVT11LL_CKT W=1.56u L=40.00n
XX13 pm CK hnet12 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX18 s CK VSS VPW NHVT11LL_CKT W=0.26u L=40.00n
XX11 cn CK VSS VPW NHVT11LL_CKT W=170.00n L=40.00n
XX17 s pm VSS VPW NHVT11LL_CKT W=0.26u L=40.00n
XX21 hnet22 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
.ENDS CLKLAHQV12_12TH40
.SUBCKT CLKLAHQV16_12TH40 CK E Q TE VDD VSS
XX6 hnet31 pm VDD VNW PHVT11LL_CKT W=1.44u L=40.00n
XX7 s CK hnet31 VNW PHVT11LL_CKT W=1.44u L=40.00n
XX9 hnet21 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX2 hnet13 TE VDD VNW PHVT11LL_CKT W=0.94u L=40.00n
XX3 hnet11 E hnet13 VNW PHVT11LL_CKT W=0.94u L=40.00n
XX5 m pm VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX10 pm CK hnet21 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 Q s VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX4 pm cn hnet11 VNW PHVT11LL_CKT W=0.94u L=40.00n
XX0 cn CK VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX20 pm cn hnet22 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 hnet12 TE VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX15 hnet12 E VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX16 m pm VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX19 Q s VSS VPW NHVT11LL_CKT W=2.08u L=40.00n
XX13 pm CK hnet12 VPW NHVT11LL_CKT W=0.47u L=40.00n
XX18 s CK VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX11 cn CK VSS VPW NHVT11LL_CKT W=170.00n L=40.00n
XX17 s pm VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX21 hnet22 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
.ENDS CLKLAHQV16_12TH40
.SUBCKT CLKLAHQV1_12TH40 CK E Q TE VDD VSS
XX6 hnet31 pm VDD VNW PHVT11LL_CKT W=0.59u L=40.00n
XX7 s CK hnet31 VNW PHVT11LL_CKT W=0.59u L=40.00n
XX9 hnet21 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX2 hnet13 TE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX3 hnet11 E hnet13 VNW PHVT11LL_CKT W=0.395u L=40.00n
XX5 m pm VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX10 pm CK hnet21 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 Q s VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX4 pm cn hnet11 VNW PHVT11LL_CKT W=0.395u L=40.00n
XX0 cn CK VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX20 pm cn hnet22 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 hnet12 TE VSS VPW NHVT11LL_CKT W=200.00n L=40.00n
XX15 hnet12 E VSS VPW NHVT11LL_CKT W=200.00n L=40.00n
XX16 m pm VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX19 Q s VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX13 pm CK hnet12 VPW NHVT11LL_CKT W=200.00n L=40.00n
XX18 s CK VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX11 cn CK VSS VPW NHVT11LL_CKT W=170.00n L=40.00n
XX17 s pm VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX21 hnet22 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
.ENDS CLKLAHQV1_12TH40
.SUBCKT CLKLAHQV20_12TH40 CK E Q TE VDD VSS
XX6 hnet31 pm VDD VNW PHVT11LL_CKT W=1.65u L=40.00n
XX7 s CK hnet31 VNW PHVT11LL_CKT W=1.65u L=40.00n
XX9 hnet21 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX2 hnet13 TE VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX3 hnet11 E hnet13 VNW PHVT11LL_CKT W=1.08u L=40.00n
XX5 m pm VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX10 pm CK hnet21 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 Q s VDD VNW PHVT11LL_CKT W=6.1u L=40.00n
XX4 pm cn hnet11 VNW PHVT11LL_CKT W=1.08u L=40.00n
XX0 cn CK VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX20 pm cn hnet22 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 hnet12 TE VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX15 hnet12 E VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX16 m pm VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX19 Q s VSS VPW NHVT11LL_CKT W=2.6u L=40.00n
XX13 pm CK hnet12 VPW NHVT11LL_CKT W=0.54u L=40.00n
XX18 s CK VSS VPW NHVT11LL_CKT W=0.39u L=40.00n
XX11 cn CK VSS VPW NHVT11LL_CKT W=170.00n L=40.00n
XX17 s pm VSS VPW NHVT11LL_CKT W=0.39u L=40.00n
XX21 hnet22 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
.ENDS CLKLAHQV20_12TH40
.SUBCKT CLKLAHQV24_12TH40 CK E Q TE VDD VSS
XX20 pm cn hnet22 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 hnet12 TE VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX15 hnet12 E VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX16 m pm VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX19 Q s VSS VPW NHVT11LL_CKT W=3.36u L=40.00n
XX13 pm CK hnet12 VPW NHVT11LL_CKT W=0.61u L=40.00n
XX18 s CK VSS VPW NHVT11LL_CKT W=0.41u L=40.00n
XX11 cn CK VSS VPW NHVT11LL_CKT W=170.00n L=40.00n
XX17 s pm VSS VPW NHVT11LL_CKT W=0.41u L=40.00n
XX21 hnet22 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX8 Q s VDD VNW PHVT11LL_CKT W=7.32u L=40.00n
XX4 pm cn hnet11 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 cn CK VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX6 hnet31 pm VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX7 s CK hnet31 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX9 hnet21 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX2 hnet13 TE VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX3 hnet11 E hnet13 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX5 m pm VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX10 pm CK hnet21 VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS CLKLAHQV24_12TH40
.SUBCKT CLKLAHQV2_12TH40 CK E Q TE VDD VSS
XX6 hnet31 pm VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX7 s CK hnet31 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX9 hnet21 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX2 hnet13 TE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX3 hnet11 E hnet13 VNW PHVT11LL_CKT W=0.44u L=40.00n
XX5 m pm VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX10 pm CK hnet21 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 Q s VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX4 pm cn hnet11 VNW PHVT11LL_CKT W=0.44u L=40.00n
XX0 cn CK VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX20 pm cn hnet22 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 hnet12 TE VSS VPW NHVT11LL_CKT W=0.22u L=40.00n
XX15 hnet12 E VSS VPW NHVT11LL_CKT W=0.22u L=40.00n
XX16 m pm VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX19 Q s VSS VPW NHVT11LL_CKT W=0.26u L=40.00n
XX13 pm CK hnet12 VPW NHVT11LL_CKT W=0.22u L=40.00n
XX18 s CK VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX11 cn CK VSS VPW NHVT11LL_CKT W=170.00n L=40.00n
XX17 s pm VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX21 hnet22 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
.ENDS CLKLAHQV2_12TH40
.SUBCKT CLKLAHQV3_12TH40 CK E Q TE VDD VSS
XX6 hnet31 pm VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX7 s CK hnet31 VNW PHVT11LL_CKT W=0.86u L=40.00n
XX9 hnet21 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX2 hnet13 TE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX3 hnet11 E hnet13 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX5 m pm VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX10 pm CK hnet21 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 Q s VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX4 pm cn hnet11 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX0 cn CK VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX20 pm cn hnet22 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 hnet12 TE VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX15 hnet12 E VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX16 m pm VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX19 Q s VSS VPW NHVT11LL_CKT W=0.37u L=40.00n
XX13 pm CK hnet12 VPW NHVT11LL_CKT W=0.23u L=40.00n
XX18 s CK VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX11 cn CK VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX17 s pm VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX21 hnet22 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
.ENDS CLKLAHQV3_12TH40
.SUBCKT CLKLAHQV4_12TH40 CK E Q TE VDD VSS
XX6 hnet31 pm VDD VNW PHVT11LL_CKT W=0.9u L=40.00n
XX7 s CK hnet31 VNW PHVT11LL_CKT W=0.9u L=40.00n
XX9 hnet21 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX2 hnet13 TE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX3 hnet11 E hnet13 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX5 m pm VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX10 pm CK hnet21 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 Q s VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX4 pm cn hnet11 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX0 cn CK VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX20 pm cn hnet22 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 hnet12 TE VSS VPW NHVT11LL_CKT W=0.24u L=40.00n
XX15 hnet12 E VSS VPW NHVT11LL_CKT W=0.24u L=40.00n
XX16 m pm VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX19 Q s VSS VPW NHVT11LL_CKT W=0.52u L=40.00n
XX13 pm CK hnet12 VPW NHVT11LL_CKT W=0.24u L=40.00n
XX18 s CK VSS VPW NHVT11LL_CKT W=0.22u L=40.00n
XX11 cn CK VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX17 s pm VSS VPW NHVT11LL_CKT W=0.22u L=40.00n
XX21 hnet22 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
.ENDS CLKLAHQV4_12TH40
.SUBCKT CLKLAHQV6_12TH40 CK E Q TE VDD VSS
XX6 hnet31 pm VDD VNW PHVT11LL_CKT W=0.9u L=40.00n
XX7 s CK hnet31 VNW PHVT11LL_CKT W=0.9u L=40.00n
XX9 hnet21 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX2 hnet13 TE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX3 hnet11 E hnet13 VNW PHVT11LL_CKT W=0.52u L=40.00n
XX5 m pm VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX10 pm CK hnet21 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 Q s VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX4 pm cn hnet11 VNW PHVT11LL_CKT W=0.52u L=40.00n
XX0 cn CK VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX20 pm cn hnet22 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 hnet12 TE VSS VPW NHVT11LL_CKT W=0.26u L=40.00n
XX15 hnet12 E VSS VPW NHVT11LL_CKT W=0.26u L=40.00n
XX16 m pm VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX19 Q s VSS VPW NHVT11LL_CKT W=0.78u L=40.00n
XX13 pm CK hnet12 VPW NHVT11LL_CKT W=0.26u L=40.00n
XX18 s CK VSS VPW NHVT11LL_CKT W=0.22u L=40.00n
XX11 cn CK VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX17 s pm VSS VPW NHVT11LL_CKT W=0.22u L=40.00n
XX21 hnet22 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
.ENDS CLKLAHQV6_12TH40
.SUBCKT CLKLAHQV8_12TH40 CK E Q TE VDD VSS
XX6 hnet31 pm VDD VNW PHVT11LL_CKT W=900.00n L=40.00n
XX7 s CK hnet31 VNW PHVT11LL_CKT W=900.00n L=40.00n
XX9 hnet21 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX2 hnet13 TE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX3 hnet11 E hnet13 VNW PHVT11LL_CKT W=0.56u L=40.00n
XX5 m pm VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX10 pm CK hnet21 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 Q s VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX4 pm cn hnet11 VNW PHVT11LL_CKT W=0.56u L=40.00n
XX0 cn CK VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX20 pm cn hnet22 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 hnet12 TE VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX15 hnet12 E VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX16 m pm VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX19 Q s VSS VPW NHVT11LL_CKT W=1.04u L=40.00n
XX13 pm CK hnet12 VPW NHVT11LL_CKT W=0.28u L=40.00n
XX18 s CK VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX11 cn CK VSS VPW NHVT11LL_CKT W=170.00n L=40.00n
XX17 s pm VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX21 hnet22 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
.ENDS CLKLAHQV8_12TH40
.SUBCKT CLKLANAQV0_12TH40 CK E Q TE VDD VSS
XX15 m pm VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
XX18 s m nt21 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX14 pm CK nt11 VNW PHVT11LL_CKT W=0.34u L=40.00n
XX13 nt11 E VDD VNW PHVT11LL_CKT W=0.34u L=40.00n
XX16 nt21 TE VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX19 Q s VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
XX20 nt13 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX17 s CK VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX21 pm cn nt13 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX3 nt12 E VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX10 nt14 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 pm cn nt12 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX0 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX4 m pm VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX8 Q s VSS VPW NHVT11LL_CKT W=130.00n L=40.00n
XX9 pm CK nt14 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 nt22 m VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX7 nt22 TE VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX5 s CK nt22 VPW NHVT11LL_CKT W=0.16u L=40.00n
.ENDS CLKLANAQV0_12TH40
.SUBCKT CLKLANAQV10_12TH40 CK E Q TE VDD VSS
XX15 m pm VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX18 s m nt21 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX14 pm CK nt11 VNW PHVT11LL_CKT W=360.00n L=40.00n
XX13 nt11 E VDD VNW PHVT11LL_CKT W=360.00n L=40.00n
XX16 nt21 TE VDD VNW PHVT11LL_CKT W=0.49u L=40.00n
XX19 Q s VDD VNW PHVT11LL_CKT W=3.05u L=40.00n
XX20 nt13 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX17 s CK VDD VNW PHVT11LL_CKT W=0.98u L=40.00n
XX21 pm cn nt13 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX3 nt12 E VSS VPW NHVT11LL_CKT W=360.00n L=40.00n
XX10 nt14 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 pm cn nt12 VPW NHVT11LL_CKT W=360.00n L=40.00n
XX0 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX4 m pm VSS VPW NHVT11LL_CKT W=0.36u L=40.00n
XX8 Q s VSS VPW NHVT11LL_CKT W=1.305u L=40.00n
XX9 pm CK nt14 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 nt22 m VSS VPW NHVT11LL_CKT W=840.00n L=40.00n
XX7 nt22 TE VSS VPW NHVT11LL_CKT W=840.00n L=40.00n
XX5 s CK nt22 VPW NHVT11LL_CKT W=840.00n L=40.00n
.ENDS CLKLANAQV10_12TH40
.SUBCKT CLKLANAQV12_12TH40 CK E Q TE VDD VSS
XX15 m pm VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX18 s m nt21 VNW PHVT11LL_CKT W=0.4u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX14 pm CK nt11 VNW PHVT11LL_CKT W=360.00n L=40.00n
XX13 nt11 E VDD VNW PHVT11LL_CKT W=360.00n L=40.00n
XX16 nt21 TE VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX19 Q s VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX20 nt13 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX17 s CK VDD VNW PHVT11LL_CKT W=1.14u L=40.00n
XX21 pm cn nt13 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX3 nt12 E VSS VPW NHVT11LL_CKT W=360.00n L=40.00n
XX10 nt14 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 pm cn nt12 VPW NHVT11LL_CKT W=360.00n L=40.00n
XX0 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX4 m pm VSS VPW NHVT11LL_CKT W=0.42u L=40.00n
XX8 Q s VSS VPW NHVT11LL_CKT W=1.56u L=40.00n
XX9 pm CK nt14 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 nt22 m VSS VPW NHVT11LL_CKT W=960.00n L=40.00n
XX7 nt22 TE VSS VPW NHVT11LL_CKT W=960.00n L=40.00n
XX5 s CK nt22 VPW NHVT11LL_CKT W=960.00n L=40.00n
.ENDS CLKLANAQV12_12TH40
.SUBCKT CLKLANAQV16_12TH40 CK E Q TE VDD VSS
XX15 m pm VDD VNW PHVT11LL_CKT W=0.48u L=40.00n
XX18 s m nt21 VNW PHVT11LL_CKT W=0.45u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX14 pm CK nt11 VNW PHVT11LL_CKT W=360.00n L=40.00n
XX13 nt11 E VDD VNW PHVT11LL_CKT W=360.00n L=40.00n
XX16 nt21 TE VDD VNW PHVT11LL_CKT W=0.45u L=40.00n
XX19 Q s VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX20 nt13 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX17 s CK VDD VNW PHVT11LL_CKT W=1.35u L=40.00n
XX21 pm cn nt13 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX3 nt12 E VSS VPW NHVT11LL_CKT W=360.00n L=40.00n
XX10 nt14 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 pm cn nt12 VPW NHVT11LL_CKT W=360.00n L=40.00n
XX0 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX4 m pm VSS VPW NHVT11LL_CKT W=0.48u L=40.00n
XX8 Q s VSS VPW NHVT11LL_CKT W=2.08u L=40.00n
XX9 pm CK nt14 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 nt22 m VSS VPW NHVT11LL_CKT W=1.17u L=40.00n
XX7 nt22 TE VSS VPW NHVT11LL_CKT W=1.17u L=40.00n
XX5 s CK nt22 VPW NHVT11LL_CKT W=1.17u L=40.00n
.ENDS CLKLANAQV16_12TH40
.SUBCKT CLKLANAQV1_12TH40 CK E Q TE VDD VSS
XX15 m pm VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
XX18 s m nt21 VNW PHVT11LL_CKT W=0.23u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX14 pm CK nt11 VNW PHVT11LL_CKT W=0.34u L=40.00n
XX13 nt11 E VDD VNW PHVT11LL_CKT W=0.34u L=40.00n
XX16 nt21 TE VDD VNW PHVT11LL_CKT W=0.23u L=40.00n
XX19 Q s VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX20 nt13 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX17 s CK VDD VNW PHVT11LL_CKT W=0.23u L=40.00n
XX21 pm cn nt13 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX3 nt12 E VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX10 nt14 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 pm cn nt12 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX0 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX4 m pm VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX8 Q s VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX9 pm CK nt14 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 nt22 m VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX7 nt22 TE VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX5 s CK nt22 VPW NHVT11LL_CKT W=0.2u L=40.00n
.ENDS CLKLANAQV1_12TH40
.SUBCKT CLKLANAQV20_12TH40 CK E Q TE VDD VSS
XX15 m pm VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX18 s m nt21 VNW PHVT11LL_CKT W=0.49u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX14 pm CK nt11 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX13 nt11 E VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
XX16 nt21 TE VDD VNW PHVT11LL_CKT W=0.49u L=40.00n
XX19 Q s VDD VNW PHVT11LL_CKT W=6.1u L=40.00n
XX20 nt13 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX17 s CK VDD VNW PHVT11LL_CKT W=1.47u L=40.00n
XX21 pm cn nt13 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX3 nt12 E VSS VPW NHVT11LL_CKT W=360.00n L=40.00n
XX10 nt14 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 pm cn nt12 VPW NHVT11LL_CKT W=360.00n L=40.00n
XX0 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX4 m pm VSS VPW NHVT11LL_CKT W=0.36u L=40.00n
XX8 Q s VSS VPW NHVT11LL_CKT W=2.6u L=40.00n
XX9 pm CK nt14 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 nt22 m VSS VPW NHVT11LL_CKT W=1.26u L=40.00n
XX7 nt22 TE VSS VPW NHVT11LL_CKT W=1.26u L=40.00n
XX5 s CK nt22 VPW NHVT11LL_CKT W=1.26u L=40.00n
.ENDS CLKLANAQV20_12TH40
.SUBCKT CLKLANAQV24_12TH40 CK E Q TE VDD VSS
XX3 nt12 E VSS VPW NHVT11LL_CKT W=360.00n L=40.00n
XX10 nt14 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 pm cn nt12 VPW NHVT11LL_CKT W=360.00n L=40.00n
XX0 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX4 m pm VSS VPW NHVT11LL_CKT W=0.6u L=40.00n
XX8 Q s VSS VPW NHVT11LL_CKT W=3.12u L=40.00n
XX9 pm CK nt14 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 nt22 m VSS VPW NHVT11LL_CKT W=1.41u L=40.00n
XX7 nt22 TE VSS VPW NHVT11LL_CKT W=1.41u L=40.00n
XX5 s CK nt22 VPW NHVT11LL_CKT W=1.41u L=40.00n
XX15 m pm VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX18 s m nt21 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX14 pm CK nt11 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX13 nt11 E VDD VNW PHVT11LL_CKT W=0.48u L=40.00n
XX16 nt21 TE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX19 Q s VDD VNW PHVT11LL_CKT W=7.32u L=40.00n
XX20 nt13 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX17 s CK VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX21 pm cn nt13 VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS CLKLANAQV24_12TH40
.SUBCKT CLKLANAQV2_12TH40 CK E Q TE VDD VSS
XX15 m pm VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
XX18 s m nt21 VNW PHVT11LL_CKT W=0.23u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX14 pm CK nt11 VNW PHVT11LL_CKT W=0.34u L=40.00n
XX13 nt11 E VDD VNW PHVT11LL_CKT W=0.34u L=40.00n
XX16 nt21 TE VDD VNW PHVT11LL_CKT W=0.23u L=40.00n
XX19 Q s VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX20 nt13 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX17 s CK VDD VNW PHVT11LL_CKT W=0.26u L=40.00n
XX21 pm cn nt13 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX3 nt12 E VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX10 nt14 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 pm cn nt12 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX0 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX4 m pm VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX8 Q s VSS VPW NHVT11LL_CKT W=0.26u L=40.00n
XX9 pm CK nt14 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 nt22 m VSS VPW NHVT11LL_CKT W=0.24u L=40.00n
XX7 nt22 TE VSS VPW NHVT11LL_CKT W=0.24u L=40.00n
XX5 s CK nt22 VPW NHVT11LL_CKT W=0.24u L=40.00n
.ENDS CLKLANAQV2_12TH40
.SUBCKT CLKLANAQV3_12TH40 CK E Q TE VDD VSS
XX15 m pm VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
XX18 s m nt21 VNW PHVT11LL_CKT W=0.24u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX14 pm CK nt11 VNW PHVT11LL_CKT W=360.00n L=40.00n
XX13 nt11 E VDD VNW PHVT11LL_CKT W=360.00n L=40.00n
XX16 nt21 TE VDD VNW PHVT11LL_CKT W=0.24u L=40.00n
XX19 Q s VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX20 nt13 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX17 s CK VDD VNW PHVT11LL_CKT W=350.00n L=40.00n
XX21 pm cn nt13 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX3 nt12 E VSS VPW NHVT11LL_CKT W=360.00n L=40.00n
XX10 nt14 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 pm cn nt12 VPW NHVT11LL_CKT W=360.00n L=40.00n
XX0 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX4 m pm VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX8 Q s VSS VPW NHVT11LL_CKT W=0.37u L=40.00n
XX9 pm CK nt14 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 nt22 m VSS VPW NHVT11LL_CKT W=280.00n L=40.00n
XX7 nt22 TE VSS VPW NHVT11LL_CKT W=280.00n L=40.00n
XX5 s CK nt22 VPW NHVT11LL_CKT W=280.00n L=40.00n
.ENDS CLKLANAQV3_12TH40
.SUBCKT CLKLANAQV4_12TH40 CK E Q TE VDD VSS
XX15 m pm VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
XX18 s m nt21 VNW PHVT11LL_CKT W=0.26u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX14 pm CK nt11 VNW PHVT11LL_CKT W=360.00n L=40.00n
XX13 nt11 E VDD VNW PHVT11LL_CKT W=360.00n L=40.00n
XX16 nt21 TE VDD VNW PHVT11LL_CKT W=0.26u L=40.00n
XX19 Q s VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX20 nt13 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX17 s CK VDD VNW PHVT11LL_CKT W=490.00n L=40.00n
XX21 pm cn nt13 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX3 nt12 E VSS VPW NHVT11LL_CKT W=360.00n L=40.00n
XX10 nt14 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 pm cn nt12 VPW NHVT11LL_CKT W=360.00n L=40.00n
XX0 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX4 m pm VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX8 Q s VSS VPW NHVT11LL_CKT W=0.52u L=40.00n
XX9 pm CK nt14 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 nt22 m VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX7 nt22 TE VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX5 s CK nt22 VPW NHVT11LL_CKT W=400.00n L=40.00n
.ENDS CLKLANAQV4_12TH40
.SUBCKT CLKLANAQV6_12TH40 CK E Q TE VDD VSS
XX15 m pm VDD VNW PHVT11LL_CKT W=0.28u L=40.00n
XX18 s m nt21 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX14 pm CK nt11 VNW PHVT11LL_CKT W=360.00n L=40.00n
XX13 nt11 E VDD VNW PHVT11LL_CKT W=360.00n L=40.00n
XX16 nt21 TE VDD VNW PHVT11LL_CKT W=0.26u L=40.00n
XX19 Q s VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX20 nt13 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX17 s CK VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX21 pm cn nt13 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX3 nt12 E VSS VPW NHVT11LL_CKT W=360.00n L=40.00n
XX10 nt14 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 pm cn nt12 VPW NHVT11LL_CKT W=360.00n L=40.00n
XX0 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX4 m pm VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX8 Q s VSS VPW NHVT11LL_CKT W=0.78u L=40.00n
XX9 pm CK nt14 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 nt22 m VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX7 nt22 TE VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX5 s CK nt22 VPW NHVT11LL_CKT W=500.00n L=40.00n
.ENDS CLKLANAQV6_12TH40
.SUBCKT CLKLANAQV8_12TH40 CK E Q TE VDD VSS
XX15 m pm VDD VNW PHVT11LL_CKT W=0.3u L=40.00n
XX18 s m nt21 VNW PHVT11LL_CKT W=0.31u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX14 pm CK nt11 VNW PHVT11LL_CKT W=360.00n L=40.00n
XX13 nt11 E VDD VNW PHVT11LL_CKT W=360.00n L=40.00n
XX16 nt21 TE VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX19 Q s VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX20 nt13 m VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX17 s CK VDD VNW PHVT11LL_CKT W=0.94u L=40.00n
XX21 pm cn nt13 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX3 nt12 E VSS VPW NHVT11LL_CKT W=360.00n L=40.00n
XX10 nt14 m VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 pm cn nt12 VPW NHVT11LL_CKT W=360.00n L=40.00n
XX0 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX4 m pm VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX8 Q s VSS VPW NHVT11LL_CKT W=1.04u L=40.00n
XX9 pm CK nt14 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 nt22 m VSS VPW NHVT11LL_CKT W=780.00n L=40.00n
XX7 nt22 TE VSS VPW NHVT11LL_CKT W=780.00n L=40.00n
XX5 s CK nt22 VPW NHVT11LL_CKT W=780.00n L=40.00n
.ENDS CLKLANAQV8_12TH40
.SUBCKT CLKLANQV0_12TH40 CK E Q TE VDD VSS
XX20 net118 TE VDD VNW PHVT11LL_CKT W=0.285u L=40.00n
XX1 net155 E net118 VNW PHVT11LL_CKT W=0.165u L=40.00n
XX3 cn CK VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX4 net155 CK net150 VNW PHVT11LL_CKT W=0.12u L=40.00n
XX6 net143 net150 VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX10 net150 cn net102 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX13 net102 net143 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX14 net127 CK VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX15 net127 net143 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX18 Q net127 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX21 net155 TE VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX2 net155 E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX0 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX5 net155 cn net150 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX7 net143 net150 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX11 net139 net143 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX12 net150 CK net139 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net131 net143 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX17 net127 CK net131 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX19 Q net127 VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
.ENDS CLKLANQV0_12TH40
.SUBCKT CLKLANQV10_12TH40 CK E Q TE VDD VSS
XX0 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX5 net87 cn net98 VPW NHVT11LL_CKT W=0.22u L=40.00n
XX21 net87 TE VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX2 net87 E VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX19 Q net115 VSS VPW NHVT11LL_CKT W=1.305u L=40.00n
XX17 net115 CK net111 VPW NHVT11LL_CKT W=0.79u L=40.00n
XX16 net111 net99 VSS VPW NHVT11LL_CKT W=0.79u L=40.00n
XX12 net98 CK net103 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX11 net103 net99 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 net99 net98 VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX18 Q net115 VDD VNW PHVT11LL_CKT W=3.05u L=40.00n
XX15 net115 net99 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX14 net115 CK VDD VNW PHVT11LL_CKT W=0.95u L=40.00n
XX13 net146 net99 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX10 net98 cn net146 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX6 net99 net98 VDD VNW PHVT11LL_CKT W=0.21u L=40.00n
XX4 net87 CK net98 VNW PHVT11LL_CKT W=0.23u L=40.00n
XX3 cn CK VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net87 E net130 VNW PHVT11LL_CKT W=0.28u L=40.00n
XX20 net130 TE VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
.ENDS CLKLANQV10_12TH40
.SUBCKT CLKLANQV12_12TH40 CK E Q TE VDD VSS
XX0 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX5 net87 cn net98 VPW NHVT11LL_CKT W=0.22u L=40.00n
XX21 net87 TE VSS VPW NHVT11LL_CKT W=0.22u L=40.00n
XX2 net87 E VSS VPW NHVT11LL_CKT W=0.22u L=40.00n
XX19 Q net115 VSS VPW NHVT11LL_CKT W=1.56u L=40.00n
XX17 net115 CK net111 VPW NHVT11LL_CKT W=0.92u L=40.00n
XX16 net111 net99 VSS VPW NHVT11LL_CKT W=0.92u L=40.00n
XX12 net98 CK net103 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX11 net103 net99 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 net99 net98 VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX18 Q net115 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX15 net115 net99 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX14 net115 CK VDD VNW PHVT11LL_CKT W=1.095u L=40.00n
XX13 net146 net99 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX10 net98 cn net146 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX6 net99 net98 VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX4 net87 CK net98 VNW PHVT11LL_CKT W=0.23u L=40.00n
XX3 cn CK VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net87 E net130 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX20 net130 TE VDD VNW PHVT11LL_CKT W=0.47u L=40.00n
.ENDS CLKLANQV12_12TH40
.SUBCKT CLKLANQV16_12TH40 CK E Q TE VDD VSS
XX0 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX5 net87 cn net98 VPW NHVT11LL_CKT W=0.265u L=40.00n
XX21 net87 TE VSS VPW NHVT11LL_CKT W=0.265u L=40.00n
XX2 net87 E VSS VPW NHVT11LL_CKT W=0.265u L=40.00n
XX19 Q net115 VSS VPW NHVT11LL_CKT W=2.08u L=40.00n
XX17 net115 CK net111 VPW NHVT11LL_CKT W=1.2u L=40.00n
XX16 net111 net99 VSS VPW NHVT11LL_CKT W=1.2u L=40.00n
XX12 net98 CK net103 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX11 net103 net99 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 net99 net98 VSS VPW NHVT11LL_CKT W=0.245u L=40.00n
XX18 Q net115 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX15 net115 net99 VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX14 net115 CK VDD VNW PHVT11LL_CKT W=1.42u L=40.00n
XX13 net146 net99 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX10 net98 cn net146 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX6 net99 net98 VDD VNW PHVT11LL_CKT W=0.28u L=40.00n
XX4 net87 CK net98 VNW PHVT11LL_CKT W=0.265u L=40.00n
XX3 cn CK VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net87 E net130 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX20 net130 TE VDD VNW PHVT11LL_CKT W=0.59u L=40.00n
.ENDS CLKLANQV16_12TH40
.SUBCKT CLKLANQV1_12TH40 CK E Q TE VDD VSS
XX0 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX5 net87 cn net98 VPW NHVT11LL_CKT W=0.16u L=40.00n
XX21 net87 TE VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX2 net87 E VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX19 Q net115 VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX17 net115 CK net111 VPW NHVT11LL_CKT W=0.16u L=40.00n
XX16 net111 net99 VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX12 net98 CK net103 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX11 net103 net99 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 net99 net98 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 Q net115 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX15 net115 net99 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX14 net115 CK VDD VNW PHVT11LL_CKT W=0.19u L=40.00n
XX13 net146 net99 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX10 net98 cn net146 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX6 net99 net98 VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX4 net87 CK net98 VNW PHVT11LL_CKT W=0.175u L=40.00n
XX3 cn CK VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net87 E net130 VNW PHVT11LL_CKT W=0.21u L=40.00n
XX20 net130 TE VDD VNW PHVT11LL_CKT W=0.37u L=40.00n
.ENDS CLKLANQV1_12TH40
.SUBCKT CLKLANQV20_12TH40 CK E Q TE VDD VSS
XX0 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX5 net87 cn net98 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX21 net87 TE VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX2 net87 E VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX19 Q net115 VSS VPW NHVT11LL_CKT W=2.6u L=40.00n
XX17 net115 CK net111 VPW NHVT11LL_CKT W=1.44u L=40.00n
XX16 net111 net99 VSS VPW NHVT11LL_CKT W=1.44u L=40.00n
XX12 net98 CK net103 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX11 net103 net99 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 net99 net98 VSS VPW NHVT11LL_CKT W=0.305u L=40.00n
XX18 Q net115 VDD VNW PHVT11LL_CKT W=6.1u L=40.00n
XX15 net115 net99 VDD VNW PHVT11LL_CKT W=0.17u L=40.00n
XX14 net115 CK VDD VNW PHVT11LL_CKT W=1.675u L=40.00n
XX13 net146 net99 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX10 net98 cn net146 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX6 net99 net98 VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX4 net87 CK net98 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX3 cn CK VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net87 E net130 VNW PHVT11LL_CKT W=0.41u L=40.00n
XX20 net130 TE VDD VNW PHVT11LL_CKT W=0.66u L=40.00n
.ENDS CLKLANQV20_12TH40
.SUBCKT CLKLANQV24_12TH40 CK E Q TE VDD VSS
XX0 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX5 net87 cn net98 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX21 net87 TE VSS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX2 net87 E VSS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX19 Q net115 VSS VPW NHVT11LL_CKT W=3.12u L=40.00n
XX17 net115 CK net111 VPW NHVT11LL_CKT W=1.68u L=40.00n
XX16 net111 net99 VSS VPW NHVT11LL_CKT W=1.68u L=40.00n
XX12 net98 CK net103 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX11 net103 net99 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 net99 net98 VSS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX18 Q net115 VDD VNW PHVT11LL_CKT W=7.32u L=40.00n
XX15 net115 net99 VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX14 net115 CK VDD VNW PHVT11LL_CKT W=1.975u L=40.00n
XX13 net146 net99 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX10 net98 cn net146 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX6 net99 net98 VDD VNW PHVT11LL_CKT W=0.375u L=40.00n
XX4 net87 CK net98 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX3 cn CK VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net87 E net130 VNW PHVT11LL_CKT W=0.45u L=40.00n
XX20 net130 TE VDD VNW PHVT11LL_CKT W=0.72u L=40.00n
.ENDS CLKLANQV24_12TH40
.SUBCKT CLKLANQV2_12TH40 CK E Q TE VDD VSS
XX0 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX5 net87 cn net98 VPW NHVT11LL_CKT W=180.00n L=40.00n
XX21 net87 TE VSS VPW NHVT11LL_CKT W=180.00n L=40.00n
XX2 net87 E VSS VPW NHVT11LL_CKT W=180.00n L=40.00n
XX19 Q net115 VSS VPW NHVT11LL_CKT W=0.26u L=40.00n
XX17 net115 CK net111 VPW NHVT11LL_CKT W=185.00n L=40.00n
XX16 net111 net99 VSS VPW NHVT11LL_CKT W=185.00n L=40.00n
XX12 net98 CK net103 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX11 net103 net99 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 net99 net98 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 Q net115 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX15 net115 net99 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX14 net115 CK VDD VNW PHVT11LL_CKT W=215.00n L=40.00n
XX13 net146 net99 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX10 net98 cn net146 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX6 net99 net98 VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX4 net87 CK net98 VNW PHVT11LL_CKT W=0.19u L=40.00n
XX3 cn CK VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net87 E net130 VNW PHVT11LL_CKT W=235.00n L=40.00n
XX20 net130 TE VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
.ENDS CLKLANQV2_12TH40
.SUBCKT CLKLANQV3_12TH40 CK E Q TE VDD VSS
XX0 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX5 net87 cn net98 VPW NHVT11LL_CKT W=0.19u L=40.00n
XX21 net87 TE VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX2 net87 E VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX19 Q net115 VSS VPW NHVT11LL_CKT W=0.37u L=40.00n
XX17 net115 CK net111 VPW NHVT11LL_CKT W=0.24u L=40.00n
XX16 net111 net99 VSS VPW NHVT11LL_CKT W=0.24u L=40.00n
XX12 net98 CK net103 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX11 net103 net99 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 net99 net98 VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX18 Q net115 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX15 net115 net99 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX14 net115 CK VDD VNW PHVT11LL_CKT W=0.29u L=40.00n
XX13 net146 net99 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX10 net98 cn net146 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX6 net99 net98 VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX4 net87 CK net98 VNW PHVT11LL_CKT W=0.19u L=40.00n
XX3 cn CK VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net87 E net130 VNW PHVT11LL_CKT W=0.25u L=40.00n
XX20 net130 TE VDD VNW PHVT11LL_CKT W=0.445u L=40.00n
.ENDS CLKLANQV3_12TH40
.SUBCKT CLKLANQV4_12TH40 CK E Q TE VDD VSS
XX0 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX5 net87 cn net98 VPW NHVT11LL_CKT W=0.19u L=40.00n
XX21 net87 TE VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX2 net87 E VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX19 Q net115 VSS VPW NHVT11LL_CKT W=0.52u L=40.00n
XX17 net115 CK net111 VPW NHVT11LL_CKT W=0.32u L=40.00n
XX16 net111 net99 VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX12 net98 CK net103 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX11 net103 net99 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 net99 net98 VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX18 Q net115 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX15 net115 net99 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX14 net115 CK VDD VNW PHVT11LL_CKT W=0.38u L=40.00n
XX13 net146 net99 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX10 net98 cn net146 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX6 net99 net98 VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX4 net87 CK net98 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX3 cn CK VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net87 E net130 VNW PHVT11LL_CKT W=0.26u L=40.00n
XX20 net130 TE VDD VNW PHVT11LL_CKT W=0.415u L=40.00n
.ENDS CLKLANQV4_12TH40
.SUBCKT CLKLANQV6_12TH40 CK E Q TE VDD VSS
XX0 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX5 net87 cn net98 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX21 net87 TE VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX2 net87 E VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX19 Q net115 VSS VPW NHVT11LL_CKT W=0.78u L=40.00n
XX17 net115 CK net111 VPW NHVT11LL_CKT W=0.46u L=40.00n
XX16 net111 net99 VSS VPW NHVT11LL_CKT W=0.46u L=40.00n
XX12 net98 CK net103 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX11 net103 net99 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 net99 net98 VSS VPW NHVT11LL_CKT W=0.145u L=40.00n
XX18 Q net115 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX15 net115 net99 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX14 net115 CK VDD VNW PHVT11LL_CKT W=0.55u L=40.00n
XX13 net146 net99 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX10 net98 cn net146 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX6 net99 net98 VDD VNW PHVT11LL_CKT W=0.165u L=40.00n
XX4 net87 CK net98 VNW PHVT11LL_CKT W=0.21u L=40.00n
XX3 cn CK VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net87 E net130 VNW PHVT11LL_CKT W=0.27u L=40.00n
XX20 net130 TE VDD VNW PHVT11LL_CKT W=0.435u L=40.00n
.ENDS CLKLANQV6_12TH40
.SUBCKT CLKLANQV8_12TH40 CK E Q TE VDD VSS
XX0 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX5 net87 cn net98 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX21 net87 TE VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX2 net87 E VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX19 Q net115 VSS VPW NHVT11LL_CKT W=1.035u L=40.00n
XX17 net115 CK net111 VPW NHVT11LL_CKT W=0.65u L=40.00n
XX16 net111 net99 VSS VPW NHVT11LL_CKT W=0.65u L=40.00n
XX12 net98 CK net103 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX11 net103 net99 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 net99 net98 VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX18 Q net115 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX15 net115 net99 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX14 net115 CK VDD VNW PHVT11LL_CKT W=0.76u L=40.00n
XX13 net146 net99 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX10 net98 cn net146 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX6 net99 net98 VDD VNW PHVT11LL_CKT W=0.185u L=40.00n
XX4 net87 CK net98 VNW PHVT11LL_CKT W=0.21u L=40.00n
XX3 cn CK VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net87 E net130 VNW PHVT11LL_CKT W=0.27u L=40.00n
XX20 net130 TE VDD VNW PHVT11LL_CKT W=0.435u L=40.00n
.ENDS CLKLANQV8_12TH40
.SUBCKT CLKMUX2V0_12TH40 I0 I1 S Z VDD VSS
XX10 SN S VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX8 Z net20 VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX5 AN SN net20 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX7 BN S net20 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX11 SN S VDD VNW PHVT11LL_CKT W=0.13u L=40.00n
XX9 Z net20 VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX4 AN S net20 VNW PHVT11LL_CKT W=0.31u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX6 BN SN net20 VNW PHVT11LL_CKT W=0.31u L=40.00n
.ENDS CLKMUX2V0_12TH40
.SUBCKT CLKMUX2V12_12TH40 I0 I1 S Z VDD VSS
XX10 SN S VSS VPW NHVT11LL_CKT W=0.73u L=40.00n
XX8 Z net20 VSS VPW NHVT11LL_CKT W=1.56u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=0.78u L=40.00n
XX5 AN SN net20 VPW NHVT11LL_CKT W=0.78u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=0.66u L=40.00n
XX7 BN S net20 VPW NHVT11LL_CKT W=0.78u L=40.00n
XX11 SN S VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX9 Z net20 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX4 AN S net20 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX6 BN SN net20 VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS CLKMUX2V12_12TH40
.SUBCKT CLKMUX2V1_12TH40 I0 I1 S Z VDD VSS
XX10 SN S VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX8 Z net20 VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX5 AN SN net20 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX7 BN S net20 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX11 SN S VDD VNW PHVT11LL_CKT W=0.13u L=40.00n
XX9 Z net20 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX4 AN S net20 VNW PHVT11LL_CKT W=0.31u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX6 BN SN net20 VNW PHVT11LL_CKT W=0.31u L=40.00n
.ENDS CLKMUX2V1_12TH40
.SUBCKT CLKMUX2V2_12TH40 I0 I1 S Z VDD VSS
XX10 SN S VSS VPW NHVT11LL_CKT W=185.00n L=40.00n
XX8 Z net20 VSS VPW NHVT11LL_CKT W=260.00n L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=185.00n L=40.00n
XX5 AN SN net20 VPW NHVT11LL_CKT W=185.00n L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=185.00n L=40.00n
XX7 BN S net20 VPW NHVT11LL_CKT W=185.00n L=40.00n
XX11 SN S VDD VNW PHVT11LL_CKT W=185.00n L=40.00n
XX9 Z net20 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX4 AN S net20 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX6 BN SN net20 VNW PHVT11LL_CKT W=430.00n L=40.00n
.ENDS CLKMUX2V2_12TH40
.SUBCKT CLKMUX2V3_12TH40 I0 I1 S Z VDD VSS
XX10 SN S VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX8 Z net20 VSS VPW NHVT11LL_CKT W=0.37u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX5 AN SN net20 VPW NHVT11LL_CKT W=0.185u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX7 BN S net20 VPW NHVT11LL_CKT W=0.185u L=40.00n
XX11 SN S VDD VNW PHVT11LL_CKT W=0.185u L=40.00n
XX9 Z net20 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX4 AN S net20 VNW PHVT11LL_CKT W=0.47u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=0.47u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=0.47u L=40.00n
XX6 BN SN net20 VNW PHVT11LL_CKT W=0.47u L=40.00n
.ENDS CLKMUX2V3_12TH40
.SUBCKT CLKMUX2V4_12TH40 I0 I1 S Z VDD VSS
XX10 SN S VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX8 Z net20 VSS VPW NHVT11LL_CKT W=0.52u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX5 AN SN net20 VPW NHVT11LL_CKT W=0.23u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX7 BN S net20 VPW NHVT11LL_CKT W=0.23u L=40.00n
XX11 SN S VDD VNW PHVT11LL_CKT W=0.23u L=40.00n
XX9 Z net20 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX4 AN S net20 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX6 BN SN net20 VNW PHVT11LL_CKT W=0.61u L=40.00n
.ENDS CLKMUX2V4_12TH40
.SUBCKT CLKMUX2V6_12TH40 I0 I1 S Z VDD VSS
XX10 SN S VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX8 Z net20 VSS VPW NHVT11LL_CKT W=0.78u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=0.37u L=40.00n
XX5 AN SN net20 VPW NHVT11LL_CKT W=0.37u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=0.37u L=40.00n
XX7 BN S net20 VPW NHVT11LL_CKT W=0.37u L=40.00n
XX11 SN S VDD VNW PHVT11LL_CKT W=0.32u L=40.00n
XX9 Z net20 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX4 AN S net20 VNW PHVT11LL_CKT W=0.86u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=1u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=0.84u L=40.00n
XX6 BN SN net20 VNW PHVT11LL_CKT W=0.86u L=40.00n
.ENDS CLKMUX2V6_12TH40
.SUBCKT CLKMUX2V8_12TH40 I0 I1 S Z VDD VSS
XX10 SN S VSS VPW NHVT11LL_CKT W=0.51u L=40.00n
XX8 Z net20 VSS VPW NHVT11LL_CKT W=1.04u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=0.48u L=40.00n
XX5 AN SN net20 VPW NHVT11LL_CKT W=0.48u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=0.44u L=40.00n
XX7 BN S net20 VPW NHVT11LL_CKT W=0.48u L=40.00n
XX11 SN S VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX9 Z net20 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX4 AN S net20 VNW PHVT11LL_CKT W=1.12u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=1.16u L=40.00n
XX6 BN SN net20 VNW PHVT11LL_CKT W=1.12u L=40.00n
.ENDS CLKMUX2V8_12TH40
.SUBCKT CLKNAND2V0_12TH40 A1 A2 ZN VDD VSS
XX2 ZN A1 net8 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX5 net8 A2 VSS VPW NHVT11LL_CKT W=260.00n L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
XX4 ZN A2 VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
.ENDS CLKNAND2V0_12TH40
.SUBCKT CLKNAND2V12_12TH40 A1 A2 ZN VDD VSS
XX2 ZN A1 net8 VPW NHVT11LL_CKT W=3.06u L=40.00n
XX5 net8 A2 VSS VPW NHVT11LL_CKT W=3.06u L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX4 ZN A2 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
.ENDS CLKNAND2V12_12TH40
.SUBCKT CLKNAND2V16_12TH40 A1 A2 ZN VDD VSS
XX2 ZN A1 net8 VPW NHVT11LL_CKT W=4.08u L=40.00n
XX5 net8 A2 VSS VPW NHVT11LL_CKT W=4.08u L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX4 ZN A2 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
.ENDS CLKNAND2V16_12TH40
.SUBCKT CLKNAND2V1_12TH40 A1 A2 ZN VDD VSS
XX2 ZN A1 net8 VPW NHVT11LL_CKT W=360.00n L=40.00n
XX5 net8 A2 VSS VPW NHVT11LL_CKT W=360.00n L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX4 ZN A2 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
.ENDS CLKNAND2V1_12TH40
.SUBCKT CLKNAND2V2_12TH40 A1 A2 ZN VDD VSS
XX2 ZN A1 net8 VPW NHVT11LL_CKT W=510.00n L=40.00n
XX5 net8 A2 VSS VPW NHVT11LL_CKT W=510.00n L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX4 ZN A2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS CLKNAND2V2_12TH40
.SUBCKT CLKNAND2V3_12TH40 A1 A2 ZN VDD VSS
XX2 ZN A1 net8 VPW NHVT11LL_CKT W=720.00n L=40.00n
XX5 net8 A2 VSS VPW NHVT11LL_CKT W=720.00n L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX4 ZN A2 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
.ENDS CLKNAND2V3_12TH40
.SUBCKT CLKNAND2V4_12TH40 A1 A2 ZN VDD VSS
XX2 ZN A1 net8 VPW NHVT11LL_CKT W=1.02u L=40.00n
XX5 net8 A2 VSS VPW NHVT11LL_CKT W=1.02u L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX4 ZN A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS CLKNAND2V4_12TH40
.SUBCKT CLKNAND2V6_12TH40 A1 A2 ZN VDD VSS
XX2 ZN A1 net8 VPW NHVT11LL_CKT W=1.53u L=40.00n
XX5 net8 A2 VSS VPW NHVT11LL_CKT W=1.53u L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX4 ZN A2 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS CLKNAND2V6_12TH40
.SUBCKT CLKNAND2V8_12TH40 A1 A2 ZN VDD VSS
XX2 ZN A1 net8 VPW NHVT11LL_CKT W=2.04u L=40.00n
XX5 net8 A2 VSS VPW NHVT11LL_CKT W=2.04u L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX4 ZN A2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS CLKNAND2V8_12TH40
.SUBCKT CLKXOR2V1_12TH40 A1 A2 Z VDD VSS
XX7 A1N A1 VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX8 net69 A1N net80 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX0 Z net80 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX4 net65 A2 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX11 net65 A1 net80 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX2 net69 net65 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX6 A1N A1 VSS VPW NHVT11LL_CKT W=185.000n L=40.00n
XX10 net65 A1N net80 VPW NHVT11LL_CKT W=185.000n L=40.00n
XX1 Z net80 VSS VPW NHVT11LL_CKT W=185.000n L=40.00n
XX3 net69 net65 VSS VPW NHVT11LL_CKT W=185.000n L=40.00n
XX5 net65 A2 VSS VPW NHVT11LL_CKT W=185.000n L=40.00n
XX9 net69 A1 net80 VPW NHVT11LL_CKT W=185.000n L=40.00n
.ENDS CLKXOR2V1_12TH40
.SUBCKT CLKXOR2V2_12TH40 A1 A2 Z VDD VSS
XX3 net57 net37 VSS VPW NHVT11LL_CKT W=260.00n L=40.00n
XX1 Z net44 VSS VPW NHVT11LL_CKT W=260.00n L=40.00n
XX6 A1N A1 VSS VPW NHVT11LL_CKT W=260.00n L=40.00n
XX9 net57 A1 net44 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX10 net37 A1N net44 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX5 net37 A2 VSS VPW NHVT11LL_CKT W=260.00n L=40.00n
XX2 net57 net37 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX0 Z net44 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX7 A1N A1 VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX8 net57 A1N net44 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX11 net37 A1 net44 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX4 net37 A2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS CLKXOR2V2_12TH40
.SUBCKT CLKXOR2V4_12TH40 A1 A2 Z VDD VSS
XX7 A1N A1 VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX8 net69 A1N net80 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX0 Z net80 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX4 net65 A2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX11 net65 A1 net80 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX2 net69 net65 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX6 A1N A1 VSS VPW NHVT11LL_CKT W=260.00n L=40.00n
XX10 net65 A1N net80 VPW NHVT11LL_CKT W=180.00n L=40.00n
XX1 Z net80 VSS VPW NHVT11LL_CKT W=520.00n L=40.00n
XX3 net69 net65 VSS VPW NHVT11LL_CKT W=260.00n L=40.00n
XX5 net65 A2 VSS VPW NHVT11LL_CKT W=260.00n L=40.00n
XX9 net69 A1 net80 VPW NHVT11LL_CKT W=180.00n L=40.00n
.ENDS CLKXOR2V4_12TH40
.SUBCKT CLKXOR2V8_12TH40 A1 A2 Z VDD VSS
XX7 A1N A1 VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX8 net69 A1N net80 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 Z net80 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX4 net65 A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX11 net65 A1 net80 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX2 net69 net65 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX6 A1N A1 VSS VPW NHVT11LL_CKT W=260.00n L=40.00n
XX10 net65 A1N net80 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX1 Z net80 VSS VPW NHVT11LL_CKT W=1.04u L=40.00n
XX3 net69 net65 VSS VPW NHVT11LL_CKT W=520.00n L=40.00n
XX5 net65 A2 VSS VPW NHVT11LL_CKT W=520.00n L=40.00n
XX9 net69 A1 net80 VPW NHVT11LL_CKT W=400.00n L=40.00n
.ENDS CLKXOR2V8_12TH40
.SUBCKT DEL2V0_12TH40 I Z VDD VSS
XX5 net2 I VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX0 Z net10 VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX2 net10 I net2 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net25 I VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX3 Z net10 VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX1 net10 I net25 VNW PHVT11LL_CKT W=0.31u L=40.00n
.ENDS DEL2V0_12TH40
.SUBCKT DEL2V2_12TH40 I Z VDD VSS
XX5 net2 I VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX0 Z net10 VSS VPW NHVT11LL_CKT W=0.26u L=40.00n
XX2 net10 I net2 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net25 I VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX3 Z net10 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 net10 I net25 VNW PHVT11LL_CKT W=0.31u L=40.00n
.ENDS DEL2V2_12TH40
.SUBCKT DEL2V4_12TH40 I Z VDD VSS
XX5 net2 I VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX0 Z net10 VSS VPW NHVT11LL_CKT W=0.52u L=40.00n
XX2 net10 I net2 VPW NHVT11LL_CKT W=0.19u L=40.00n
XX4 net25 I VDD VNW PHVT11LL_CKT W=0.55u L=40.00n
XX3 Z net10 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 net10 I net25 VNW PHVT11LL_CKT W=0.55u L=40.00n
.ENDS DEL2V4_12TH40
.SUBCKT DEL2V8_12TH40 I Z VDD VSS
XX5 net2 I VSS VPW NHVT11LL_CKT W=0.42u L=40.00n
XX0 Z net10 VSS VPW NHVT11LL_CKT W=1.04u L=40.00n
XX2 net10 I net2 VPW NHVT11LL_CKT W=0.42u L=40.00n
XX4 net25 I VDD VNW PHVT11LL_CKT W=0.98u L=40.00n
XX3 Z net10 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 net10 I net25 VNW PHVT11LL_CKT W=0.98u L=40.00n
.ENDS DEL2V8_12TH40
.SUBCKT DEL4V0_12TH40 I Z VDD VSS
XX13 net35 net47 net39 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX12 net39 net47 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net43 net51 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX8 net47 net51 net43 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net51 I net55 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX0 Z net35 VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX5 net55 I VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX11 net35 net47 net10 VNW PHVT11LL_CKT W=0.31u L=40.00n
XX10 net10 net47 VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX7 net22 net51 VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX6 net47 net51 net22 VNW PHVT11LL_CKT W=0.31u L=40.00n
XX1 net51 I net26 VNW PHVT11LL_CKT W=0.31u L=40.00n
XX3 Z net35 VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX4 net26 I VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
.ENDS DEL4V0_12TH40
.SUBCKT DEL4V2_12TH40 I Z VDD VSS
XX13 net35 net47 net39 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX12 net39 net47 VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX9 net43 net51 VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX8 net47 net51 net43 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX2 net51 I net55 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX0 Z net35 VSS VPW NHVT11LL_CKT W=0.26u L=40.00n
XX5 net55 I VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX11 net35 net47 net10 VNW PHVT11LL_CKT W=0.31u L=40.00n
XX10 net10 net47 VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX7 net22 net51 VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX6 net47 net51 net22 VNW PHVT11LL_CKT W=0.31u L=40.00n
XX1 net51 I net26 VNW PHVT11LL_CKT W=0.31u L=40.00n
XX3 Z net35 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX4 net26 I VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
.ENDS DEL4V2_12TH40
.SUBCKT DEL4V4_12TH40 I Z VDD VSS
XX13 net35 net47 net39 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX12 net39 net47 VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX9 net43 net51 VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX8 net47 net51 net43 VPW NHVT11LL_CKT W=0.185u L=40.00n
XX2 net51 I net55 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX0 Z net35 VSS VPW NHVT11LL_CKT W=0.52u L=40.00n
XX5 net55 I VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX11 net35 net47 net10 VNW PHVT11LL_CKT W=0.425u L=40.00n
XX10 net10 net47 VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX7 net22 net51 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX6 net47 net51 net22 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX1 net51 I net26 VNW PHVT11LL_CKT W=0.31u L=40.00n
XX3 Z net35 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX4 net26 I VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
.ENDS DEL4V4_12TH40
.SUBCKT DEL4V8_12TH40 I Z VDD VSS
XX13 net35 net47 net39 VPW NHVT11LL_CKT W=0.37u L=40.00n
XX12 net39 net47 VSS VPW NHVT11LL_CKT W=0.37u L=40.00n
XX9 net43 net51 VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX8 net47 net51 net43 VPW NHVT11LL_CKT W=0.185u L=40.00n
XX2 net51 I net55 VPW NHVT11LL_CKT W=0.185u L=40.00n
XX0 Z net35 VSS VPW NHVT11LL_CKT W=1.04u L=40.00n
XX5 net55 I VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX11 net35 net47 net10 VNW PHVT11LL_CKT W=0.86u L=40.00n
XX10 net10 net47 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX7 net22 net51 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX6 net47 net51 net22 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX1 net51 I net26 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX3 Z net35 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX4 net26 I VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
.ENDS DEL4V8_12TH40
.SUBCKT DGRNQNV2_12TH40 CK D QN RN VDD VSS
XX27 net_5 cn pm VPW NHVT11LL_CKT W=0.4u L=40.00n
XX25 QN net43 VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX1 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX4 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX8 net_5 D net_61 VPW NHVT11LL_CKT W=0.5u L=40.00n
XX9 net_61 RN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX11 m pm VSS VPW NHVT11LL_CKT W=0.475u L=40.00n
XX19 net_85 net43 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX17 m c net43 VPW NHVT11LL_CKT W=0.39u L=40.00n
XX14 net_100 c pm VPW NHVT11LL_CKT W=120.00n L=40.00n
XX15 VSS m net_100 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 net_108 cn net43 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX23 VSS net_85 net_108 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net_5 c pm VNW PHVT11LL_CKT W=0.33u L=40.00n
XX24 QN net43 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX2 net_5 RN VDD VNW PHVT11LL_CKT W=0.27u L=40.00n
XX3 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX10 m pm VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX12 VDD m net_53 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX16 m cn net43 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX18 net_85 net43 VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX20 VDD net_85 net_49 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX21 net_49 c net43 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX13 net_53 cn pm VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net_5 D VDD VNW PHVT11LL_CKT W=0.27u L=40.00n
.ENDS DGRNQNV2_12TH40
.SUBCKT DGRNQNV4_12TH40 CK D QN RN VDD VSS
XX27 net_5 cn pm VPW NHVT11LL_CKT W=0.43u L=40.00n
XX25 QN net43 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX1 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX4 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX8 net_5 D net_61 VPW NHVT11LL_CKT W=0.53u L=40.00n
XX9 net_61 RN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX11 m pm VSS VPW NHVT11LL_CKT W=0.475u L=40.00n
XX19 net_85 net43 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX17 m c net43 VPW NHVT11LL_CKT W=0.39u L=40.00n
XX14 net_100 c pm VPW NHVT11LL_CKT W=120.00n L=40.00n
XX15 VSS m net_100 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 net_108 cn net43 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX23 VSS net_85 net_108 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net_5 c pm VNW PHVT11LL_CKT W=0.33u L=40.00n
XX24 QN net43 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX2 net_5 RN VDD VNW PHVT11LL_CKT W=0.27u L=40.00n
XX3 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX10 m pm VDD VNW PHVT11LL_CKT W=0.55u L=40.00n
XX12 VDD m net_53 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX16 m cn net43 VNW PHVT11LL_CKT W=0.4u L=40.00n
XX18 net_85 net43 VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX20 VDD net_85 net_49 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX21 net_49 c net43 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX13 net_53 cn pm VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net_5 D VDD VNW PHVT11LL_CKT W=0.27u L=40.00n
.ENDS DGRNQNV4_12TH40
.SUBCKT DGRNQNV6_12TH40 CK D QN RN VDD VSS
XX27 net_5 cn pm VPW NHVT11LL_CKT W=0.335u L=40.00n
XX25 QN net43 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX1 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX4 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX8 net_5 D net_61 VPW NHVT11LL_CKT W=0.61u L=40.00n
XX9 net_61 RN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX11 m pm VSS VPW NHVT11LL_CKT W=0.435u L=40.00n
XX19 net_85 net43 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX17 m c net43 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX14 net_100 c pm VPW NHVT11LL_CKT W=120.00n L=40.00n
XX15 VSS m net_100 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 net_108 cn net43 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX23 VSS net_85 net_108 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net_5 c pm VNW PHVT11LL_CKT W=0.33u L=40.00n
XX24 QN net43 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX0 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX2 net_5 RN VDD VNW PHVT11LL_CKT W=0.3u L=40.00n
XX3 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX10 m pm VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX12 VDD m net_53 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX16 m cn net43 VNW PHVT11LL_CKT W=0.45u L=40.00n
XX18 net_85 net43 VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX20 VDD net_85 net_49 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX21 net_49 c net43 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX13 net_53 cn pm VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net_5 D VDD VNW PHVT11LL_CKT W=0.3u L=40.00n
.ENDS DGRNQNV6_12TH40
.SUBCKT DGRNQV2_12TH40 CK D Q RN VDD VSS
XX27 net_5 cn pm VPW NHVT11LL_CKT W=0.33u L=40.00n
XX25 Q net_85 VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX1 cn CK VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX4 c cn VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX8 net_5 D net_61 VPW NHVT11LL_CKT W=0.5u L=40.00n
XX9 net_61 RN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX11 m pm VSS VPW NHVT11LL_CKT W=0.415u L=40.00n
XX19 net_85 net43 VSS VPW NHVT11LL_CKT W=0.24u L=40.00n
XX17 m c net43 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX14 net_100 c pm VPW NHVT11LL_CKT W=120.00n L=40.00n
XX15 VSS m net_100 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 net_108 cn net43 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX23 VSS net_85 net_108 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net_5 c pm VNW PHVT11LL_CKT W=0.33u L=40.00n
XX24 Q net_85 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX2 net_5 RN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX3 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX10 m pm VDD VNW PHVT11LL_CKT W=0.495u L=40.00n
XX12 VDD m net_53 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX16 m cn net43 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX18 net_85 net43 VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX20 VDD net_85 net_49 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX21 net_49 c net43 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX13 net_53 cn pm VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net_5 D VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
.ENDS DGRNQV2_12TH40
.SUBCKT DGRNQV4_12TH40 CK D Q RN VDD VSS
XX27 net_5 cn pm VPW NHVT11LL_CKT W=0.33u L=40.00n
XX25 Q net_85 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX1 cn CK VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX4 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX8 net_5 D net_61 VPW NHVT11LL_CKT W=0.5u L=40.00n
XX9 net_61 RN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX11 m pm VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX19 net_85 net43 VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX17 m c net43 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX14 net_100 c pm VPW NHVT11LL_CKT W=120.00n L=40.00n
XX15 VSS m net_100 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 net_108 cn net43 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX23 VSS net_85 net_108 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net_5 c pm VNW PHVT11LL_CKT W=0.33u L=40.00n
XX24 Q net_85 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX2 net_5 RN VDD VNW PHVT11LL_CKT W=0.27u L=40.00n
XX3 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX10 m pm VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX12 VDD m net_53 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX16 m cn net43 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX18 net_85 net43 VDD VNW PHVT11LL_CKT W=0.51u L=40.00n
XX20 VDD net_85 net_49 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX21 net_49 c net43 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX13 net_53 cn pm VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net_5 D VDD VNW PHVT11LL_CKT W=0.27u L=40.00n
.ENDS DGRNQV4_12TH40
.SUBCKT DGRNQV6_12TH40 CK D Q RN VDD VSS
XX27 net_5 cn pm VPW NHVT11LL_CKT W=0.33u L=40.00n
XX25 Q net_85 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX1 cn CK VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX4 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX8 net_5 D net_61 VPW NHVT11LL_CKT W=0.61u L=40.00n
XX9 net_61 RN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX11 m pm VSS VPW NHVT11LL_CKT W=0.475u L=40.00n
XX19 net_85 net43 VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX17 m c net43 VPW NHVT11LL_CKT W=0.39u L=40.00n
XX14 net_100 c pm VPW NHVT11LL_CKT W=120.00n L=40.00n
XX15 VSS m net_100 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 net_108 cn net43 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX23 VSS net_85 net_108 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net_5 c pm VNW PHVT11LL_CKT W=0.33u L=40.00n
XX24 Q net_85 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX0 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX2 net_5 RN VDD VNW PHVT11LL_CKT W=0.3u L=40.00n
XX3 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX10 m pm VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX12 VDD m net_53 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX16 m cn net43 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX18 net_85 net43 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX20 VDD net_85 net_49 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX21 net_49 c net43 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX13 net_53 cn pm VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net_5 D VDD VNW PHVT11LL_CKT W=0.3u L=40.00n
.ENDS DGRNQV6_12TH40
.SUBCKT DGRSNQNV2_12TH40 CK D QN RN SN VDD VSS
XX30 net_66 cn net051 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX25 QN net073 VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX9 net_17 RN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX8 net_66 D net_17 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX3 net_66 snn net_17 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX13 net049 net051 VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX23 net_30 net073 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX21 net049 c net073 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX17 VSS net049 net_41 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX28 net_49 cn net073 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 VSS net_30 net_49 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 cn CK VSS VPW NHVT11LL_CKT W=130.00n L=40.00n
XX11 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX19 snn SN VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX16 net_41 c net051 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net_66 c net051 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX20 net049 cn net073 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX22 net_30 net073 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX0 net_66 RN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX24 QN net073 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX5 net_66 D net_73 VNW PHVT11LL_CKT W=0.47u L=40.00n
XX4 net_73 snn VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX12 net049 net051 VDD VNW PHVT11LL_CKT W=0.455u L=40.00n
XX14 VDD net049 net_102 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net_102 cn net051 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX26 VDD net_30 net_110 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX27 net_110 c net073 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX1 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX10 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX18 snn SN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
.ENDS DGRSNQNV2_12TH40
.SUBCKT DGRSNQNV4_12TH40 CK D QN RN SN VDD VSS
XX30 net_66 cn net051 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX25 QN net073 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX9 net_17 RN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX8 net_66 D net_17 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX3 net_66 snn net_17 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX13 net049 net051 VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX23 net_30 net073 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX21 net049 c net073 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX17 VSS net049 net_41 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX28 net_49 cn net073 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 VSS net_30 net_49 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 cn CK VSS VPW NHVT11LL_CKT W=130.00n L=40.00n
XX11 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX19 snn SN VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX16 net_41 c net051 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net_66 c net051 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX20 net049 cn net073 VNW PHVT11LL_CKT W=0.39u L=40.00n
XX22 net_30 net073 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX0 net_66 RN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX24 QN net073 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX5 net_66 D net_73 VNW PHVT11LL_CKT W=0.545u L=40.00n
XX4 net_73 snn VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX12 net049 net051 VDD VNW PHVT11LL_CKT W=0.53u L=40.00n
XX14 VDD net049 net_102 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net_102 cn net051 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX26 VDD net_30 net_110 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX27 net_110 c net073 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX1 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX10 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX18 snn SN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
.ENDS DGRSNQNV4_12TH40
.SUBCKT DGRSNQNV6_12TH40 CK D QN RN SN VDD VSS
XX30 net_66 cn net051 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX25 QN net073 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX9 net_17 RN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX8 net_66 D net_17 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX3 net_66 snn net_17 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX13 net049 net051 VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX23 net_30 net073 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX21 net049 c net073 VPW NHVT11LL_CKT W=0.37u L=40.00n
XX17 VSS net049 net_41 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX28 net_49 cn net073 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 VSS net_30 net_49 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 cn CK VSS VPW NHVT11LL_CKT W=130.00n L=40.00n
XX11 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX19 snn SN VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX16 net_41 c net051 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net_66 c net051 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX20 net049 cn net073 VNW PHVT11LL_CKT W=0.425u L=40.00n
XX22 net_30 net073 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX0 net_66 RN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX24 QN net073 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX5 net_66 D net_73 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX4 net_73 snn VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX12 net049 net051 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX14 VDD net049 net_102 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net_102 cn net051 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX26 VDD net_30 net_110 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX27 net_110 c net073 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX1 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX10 c cn VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX18 snn SN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
.ENDS DGRSNQNV6_12TH40
.SUBCKT DGRSNQV2_12TH40 CK D Q RN SN VDD VSS
XX30 net_66 cn net051 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX25 Q net_30 VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX9 net_17 RN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX8 net_66 D net_17 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX3 net_66 snn net_17 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX13 net049 net051 VSS VPW NHVT11LL_CKT W=0.45u L=40.00n
XX23 net_30 net073 VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX21 net049 c net073 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX17 VSS net049 net_41 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX28 net_49 cn net073 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 VSS net_30 net_49 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 cn CK VSS VPW NHVT11LL_CKT W=130.00n L=40.00n
XX11 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX19 snn SN VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX16 net_41 c net051 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net_66 c net051 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX20 net049 cn net073 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX22 net_30 net073 VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX0 net_66 RN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX24 Q net_30 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX5 net_66 D net_73 VNW PHVT11LL_CKT W=0.47u L=40.00n
XX4 net_73 snn VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX12 net049 net051 VDD VNW PHVT11LL_CKT W=0.45u L=40.00n
XX14 VDD net049 net_102 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net_102 cn net051 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX26 VDD net_30 net_110 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX27 net_110 c net073 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX1 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX10 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX18 snn SN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
.ENDS DGRSNQV2_12TH40
.SUBCKT DGRSNQV4_12TH40 CK D Q RN SN VDD VSS
XX30 net_66 cn net051 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX25 Q net_30 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX9 net_17 RN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX8 net_66 D net_17 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX3 net_66 snn net_17 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX13 net049 net051 VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX23 net_30 net073 VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX21 net049 c net073 VPW NHVT11LL_CKT W=0.37u L=40.00n
XX17 VSS net049 net_41 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX28 net_49 cn net073 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 VSS net_30 net_49 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 cn CK VSS VPW NHVT11LL_CKT W=130.00n L=40.00n
XX11 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX19 snn SN VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX16 net_41 c net051 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net_66 c net051 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX20 net049 cn net073 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX22 net_30 net073 VDD VNW PHVT11LL_CKT W=0.51u L=40.00n
XX0 net_66 RN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX24 Q net_30 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX5 net_66 D net_73 VNW PHVT11LL_CKT W=0.545u L=40.00n
XX4 net_73 snn VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX12 net049 net051 VDD VNW PHVT11LL_CKT W=0.495u L=40.00n
XX14 VDD net049 net_102 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net_102 cn net051 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX26 VDD net_30 net_110 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX27 net_110 c net073 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX1 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX10 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX18 snn SN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
.ENDS DGRSNQV4_12TH40
.SUBCKT DGRSNQV6_12TH40 CK D Q RN SN VDD VSS
XX30 net_66 cn net051 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX25 Q net_30 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX9 net_17 RN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX8 net_66 D net_17 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX3 net_66 snn net_17 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX13 net049 net051 VSS VPW NHVT11LL_CKT W=0.52u L=40.00n
XX23 net_30 net073 VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX21 net049 c net073 VPW NHVT11LL_CKT W=0.42u L=40.00n
XX17 VSS net049 net_41 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX28 net_49 cn net073 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 VSS net_30 net_49 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 cn CK VSS VPW NHVT11LL_CKT W=130.00n L=40.00n
XX11 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX19 snn SN VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX16 net_41 c net051 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net_66 c net051 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX20 net049 cn net073 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX22 net_30 net073 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net_66 RN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX24 Q net_30 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX5 net_66 D net_73 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX4 net_73 snn VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX12 net049 net051 VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX14 VDD net049 net_102 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net_102 cn net051 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX26 VDD net_30 net_110 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX27 net_110 c net073 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX1 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX10 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX18 snn SN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
.ENDS DGRSNQV6_12TH40
.SUBCKT DGSNQNV2_12TH40 CK D QN SN VDD VSS
XX28 net_85 cn net051 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX27 VSS net_81 net_64 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net_64 cn net073 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX15 VSS net049 net_72 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX19 net049 c net073 VPW NHVT11LL_CKT W=0.37u L=40.00n
XX11 net049 net051 VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX21 net_81 net073 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net_85 snn VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX17 snn SN VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX9 net_85 D VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX1 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX4 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX23 QN net073 VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX14 net_72 c net051 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 net_85 c net051 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX13 net_5 cn net051 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 VDD net_81 net_57 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX18 net049 cn net073 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX12 VDD net049 net_5 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX10 net049 net051 VDD VNW PHVT11LL_CKT W=0.495u L=40.00n
XX20 net_81 net073 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX6 net_85 D net_32 VNW PHVT11LL_CKT W=0.47u L=40.00n
XX5 net_32 snn VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX16 snn SN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX3 c cn VDD VNW PHVT11LL_CKT W=0.47u L=40.00n
XX0 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX22 QN net073 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX25 net_57 c net073 VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS DGSNQNV2_12TH40
.SUBCKT DGSNQNV4_12TH40 CK D QN SN VDD VSS
XX28 net_85 cn net051 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX27 VSS net_81 net_64 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net_64 cn net073 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX15 VSS net049 net_72 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX19 net049 c net073 VPW NHVT11LL_CKT W=0.37u L=40.00n
XX11 net049 net051 VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX21 net_81 net073 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net_85 snn VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX17 snn SN VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX9 net_85 D VSS VPW NHVT11LL_CKT W=0.26u L=40.00n
XX1 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX4 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX23 QN net073 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX14 net_72 c net051 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 net_85 c net051 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX13 net_5 cn net051 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 VDD net_81 net_57 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX18 net049 cn net073 VNW PHVT11LL_CKT W=0.4u L=40.00n
XX12 VDD net049 net_5 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX10 net049 net051 VDD VNW PHVT11LL_CKT W=0.55u L=40.00n
XX20 net_81 net073 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX6 net_85 D net_32 VNW PHVT11LL_CKT W=0.54u L=40.00n
XX5 net_32 snn VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX16 snn SN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX3 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX0 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX22 QN net073 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX25 net_57 c net073 VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS DGSNQNV4_12TH40
.SUBCKT DGSNQNV6_12TH40 CK D QN SN VDD VSS
XX28 net_85 cn net051 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX27 VSS net_81 net_64 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net_64 cn net073 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX15 VSS net049 net_72 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX19 net049 c net073 VPW NHVT11LL_CKT W=0.37u L=40.00n
XX11 net049 net051 VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX21 net_81 net073 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net_85 snn VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX17 snn SN VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX9 net_85 D VSS VPW NHVT11LL_CKT W=0.26u L=40.00n
XX1 cn CK VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX4 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX23 QN net073 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX14 net_72 c net051 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 net_85 c net051 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX13 net_5 cn net051 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 VDD net_81 net_57 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX18 net049 cn net073 VNW PHVT11LL_CKT W=0.425u L=40.00n
XX12 VDD net049 net_5 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX10 net049 net051 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX20 net_81 net073 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX6 net_85 D net_32 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX5 net_32 snn VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX16 snn SN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX3 c cn VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX0 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX22 QN net073 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX25 net_57 c net073 VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS DGSNQNV6_12TH40
.SUBCKT DGSNQV2_12TH40 CK D Q SN VDD VSS
XX28 net_85 cn net051 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX27 VSS net_81 net_64 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net_64 cn net073 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX15 VSS net049 net_72 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX19 net049 c net073 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX11 net049 net051 VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX21 net_81 net073 VSS VPW NHVT11LL_CKT W=0.26u L=40.00n
XX2 net_85 snn VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX17 snn SN VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX9 net_85 D VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX1 cn CK VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX4 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX23 Q net_81 VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX14 net_72 c net051 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 net_85 c net051 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX13 net_5 cn net051 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 VDD net_81 net_57 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX18 net049 cn net073 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX12 VDD net049 net_5 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX10 net049 net051 VDD VNW PHVT11LL_CKT W=0.495u L=40.00n
XX20 net_81 net073 VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX6 net_85 D net_32 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX5 net_32 snn VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX16 snn SN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX3 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX0 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX22 Q net_81 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX25 net_57 c net073 VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS DGSNQV2_12TH40
.SUBCKT DGSNQV4_12TH40 CK D Q SN VDD VSS
XX28 net_85 cn net051 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX27 VSS net_81 net_64 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net_64 cn net073 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX15 VSS net049 net_72 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX19 net049 c net073 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX11 net049 net051 VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX21 net_81 net073 VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX2 net_85 snn VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX17 snn SN VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX9 net_85 D VSS VPW NHVT11LL_CKT W=0.26u L=40.00n
XX1 cn CK VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX4 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX23 Q net_81 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX14 net_72 c net051 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 net_85 c net051 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX13 net_5 cn net051 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 VDD net_81 net_57 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX18 net049 cn net073 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX12 VDD net049 net_5 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX10 net049 net051 VDD VNW PHVT11LL_CKT W=0.495u L=40.00n
XX20 net_81 net073 VDD VNW PHVT11LL_CKT W=0.51u L=40.00n
XX6 net_85 D net_32 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX5 net_32 snn VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX16 snn SN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX3 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX0 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX22 Q net_81 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX25 net_57 c net073 VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS DGSNQV4_12TH40
.SUBCKT DGSNQV6_12TH40 CK D Q SN VDD VSS
XX28 net_85 cn net051 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX27 VSS net_81 net_64 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net_64 cn net073 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX15 VSS net049 net_72 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX19 net049 c net073 VPW NHVT11LL_CKT W=0.37u L=40.00n
XX11 net049 net051 VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX21 net_81 net073 VSS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX2 net_85 snn VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX17 snn SN VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX9 net_85 D VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX1 cn CK VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX4 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX23 Q net_81 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX14 net_72 c net051 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 net_85 c net051 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX13 net_5 cn net051 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 VDD net_81 net_57 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX18 net049 cn net073 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX12 VDD net049 net_5 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX10 net049 net051 VDD VNW PHVT11LL_CKT W=0.495u L=40.00n
XX20 net_81 net073 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX6 net_85 D net_32 VNW PHVT11LL_CKT W=0.51u L=40.00n
XX5 net_32 snn VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX16 snn SN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX3 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX0 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX22 Q net_81 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX25 net_57 c net073 VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS DGSNQV6_12TH40
.SUBCKT DQNV0_12TH40 CK D QN VDD VSS
XX2 net56 D VSS VPW NHVT11LL_CKT W=0.36u L=40.00n
XX3 net56 cn net63 VPW NHVT11LL_CKT W=0.24u L=40.00n
XX4 net64 net63 VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX6 net63 c net72 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net72 net64 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX14 net64 c net87 VPW NHVT11LL_CKT W=0.245u L=40.00n
XX16 net88 net96 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net87 cn net88 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net96 net87 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net87 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX1 net56 D VDD VNW PHVT11LL_CKT W=0.24u L=40.00n
XX0 net56 c net63 VNW PHVT11LL_CKT W=0.22u L=40.00n
XX5 net64 net63 VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX7 net63 cn net23 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net23 net64 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.13u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX15 net64 cn net87 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX19 net47 net96 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net87 c net47 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX21 net96 net87 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net87 VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
.ENDS DQNV0_12TH40
.SUBCKT DQNV2_12TH40 CK D QN VDD VSS
XX2 net56 D VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX3 net56 cn net63 VPW NHVT11LL_CKT W=330.00n L=40.00n
XX4 net64 net63 VSS VPW NHVT11LL_CKT W=0.475u L=40.00n
XX6 net63 c net72 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net72 net64 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=190.00n L=40.00n
XX14 net64 c net87 VPW NHVT11LL_CKT W=0.35u L=40.00n
XX16 net88 net96 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net87 cn net88 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net96 net87 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net87 VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX1 net56 D VDD VNW PHVT11LL_CKT W=0.26u L=40.00n
XX0 net56 c net63 VNW PHVT11LL_CKT W=0.26u L=40.00n
XX5 net64 net63 VDD VNW PHVT11LL_CKT W=0.53u L=40.00n
XX7 net63 cn net23 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net23 net64 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.13u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX15 net64 cn net87 VNW PHVT11LL_CKT W=0.31u L=40.00n
XX19 net47 net96 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net87 c net47 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX21 net96 net87 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net87 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS DQNV2_12TH40
.SUBCKT DQNV4_12TH40 CK D QN VDD VSS
XX2 net56 D VSS VPW NHVT11LL_CKT W=0.46u L=40.00n
XX3 net56 cn net63 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX4 net64 net63 VSS VPW NHVT11LL_CKT W=0.46u L=40.00n
XX6 net63 c net72 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net72 net64 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.155u L=40.00n
XX14 net64 c net87 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX16 net88 net96 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net87 cn net88 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net96 net87 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net87 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX1 net56 D VDD VNW PHVT11LL_CKT W=0.32u L=40.00n
XX0 net56 c net63 VNW PHVT11LL_CKT W=0.26u L=40.00n
XX5 net64 net63 VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX7 net63 cn net23 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net23 net64 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX15 net64 cn net87 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX19 net47 net96 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net87 c net47 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX21 net96 net87 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net87 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS DQNV4_12TH40
.SUBCKT DQNV6_12TH40 CK D QN VDD VSS
XX2 net56 D VSS VPW NHVT11LL_CKT W=0.59u L=40.00n
XX3 net56 cn net63 VPW NHVT11LL_CKT W=0.5u L=40.00n
XX4 net64 net63 VSS VPW NHVT11LL_CKT W=0.49u L=40.00n
XX6 net63 c net72 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net72 net64 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX14 net64 c net87 VPW NHVT11LL_CKT W=0.35u L=40.00n
XX16 net88 net96 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net87 cn net88 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net96 net87 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net87 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX1 net56 D VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX0 net56 c net63 VNW PHVT11LL_CKT W=0.42u L=40.00n
XX5 net64 net63 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX7 net63 cn net23 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net23 net64 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.21u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX15 net64 cn net87 VNW PHVT11LL_CKT W=0.54u L=40.00n
XX19 net47 net96 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net87 c net47 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX21 net96 net87 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net87 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS DQNV6_12TH40
.SUBCKT DQV0_12TH40 CK D Q VDD VSS
XX22 Q net8 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX18 net8 net23 VSS VPW NHVT11LL_CKT W=0.135u L=40.00n
XX17 net23 cn net16 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net16 net8 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net40 c net23 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX9 net32 net40 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net40 net47 VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX3 net48 cn net47 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX2 net48 D VSS VPW NHVT11LL_CKT W=0.305u L=40.00n
XX6 net47 c net32 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX23 Q net8 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX21 net8 net23 VDD VNW PHVT11LL_CKT W=0.24u L=40.00n
XX20 net23 c net63 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net63 net8 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net40 cn net23 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.38u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX8 net87 net40 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net47 cn net87 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net40 net47 VDD VNW PHVT11LL_CKT W=440.00n L=40.00n
XX0 net48 c net47 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX1 net48 D VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
.ENDS DQV0_12TH40
.SUBCKT DQV2_12TH40 CK D Q VDD VSS
XX22 Q net8 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX18 net8 net23 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX17 net23 cn net16 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net16 net8 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net40 c net23 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=185.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=130.00n L=40.00n
XX9 net32 net40 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net40 net47 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX3 net48 cn net47 VPW NHVT11LL_CKT W=0.28u L=40.00n
XX2 net48 D VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX6 net47 c net32 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX23 Q net8 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX21 net8 net23 VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX20 net23 c net63 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net63 net8 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net40 cn net23 VNW PHVT11LL_CKT W=0.28u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX8 net87 net40 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net47 cn net87 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net40 net47 VDD VNW PHVT11LL_CKT W=440.00n L=40.00n
XX0 net48 c net47 VNW PHVT11LL_CKT W=0.25u L=40.00n
XX1 net48 D VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
.ENDS DQV2_12TH40
.SUBCKT DQV4_12TH40 CK D Q VDD VSS
XX22 Q net8 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX18 net8 net23 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX17 net23 cn net16 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net16 net8 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net40 c net23 VPW NHVT11LL_CKT W=0.34u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX9 net32 net40 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net40 net47 VSS VPW NHVT11LL_CKT W=0.42u L=40.00n
XX3 net48 cn net47 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX2 net48 D VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX6 net47 c net32 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX23 Q net8 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX21 net8 net23 VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX20 net23 c net63 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net63 net8 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net40 cn net23 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.18u L=40.00n
XX8 net87 net40 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net47 cn net87 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net40 net47 VDD VNW PHVT11LL_CKT W=0.48u L=40.00n
XX0 net48 c net47 VNW PHVT11LL_CKT W=0.27u L=40.00n
XX1 net48 D VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
.ENDS DQV4_12TH40
.SUBCKT DQV6_12TH40 CK D Q VDD VSS
XX22 Q net8 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX18 net8 net23 VSS VPW NHVT11LL_CKT W=0.37u L=40.00n
XX17 net23 cn net16 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net16 net8 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net40 c net23 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX9 net32 net40 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net40 net47 VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX3 net48 cn net47 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX2 net48 D VSS VPW NHVT11LL_CKT W=0.48u L=40.00n
XX6 net47 c net32 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX23 Q net8 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX21 net8 net23 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX20 net23 c net63 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net63 net8 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net40 cn net23 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX8 net87 net40 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net47 cn net87 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net40 net47 VDD VNW PHVT11LL_CKT W=0.57u L=40.00n
XX0 net48 c net47 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX1 net48 D VDD VNW PHVT11LL_CKT W=0.39u L=40.00n
.ENDS DQV6_12TH40
.SUBCKT DQV8_12TH40 CK D Q VDD VSS
XX22 Q net8 VSS VPW NHVT11LL_CKT W=2.14u L=40.00n
XX18 net8 net23 VSS VPW NHVT11LL_CKT W=0.64u L=40.00n
XX17 net23 cn net16 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net16 net8 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net40 c net23 VPW NHVT11LL_CKT W=0.44u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX9 net32 net40 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net40 net47 VSS VPW NHVT11LL_CKT W=0.53u L=40.00n
XX3 net48 cn net47 VPW NHVT11LL_CKT W=0.5u L=40.00n
XX2 net48 D VSS VPW NHVT11LL_CKT W=0.59u L=40.00n
XX6 net47 c net32 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX23 Q net8 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX21 net8 net23 VDD VNW PHVT11LL_CKT W=0.88u L=40.00n
XX20 net23 c net63 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net63 net8 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net40 cn net23 VNW PHVT11LL_CKT W=0.49u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.21u L=40.00n
XX8 net87 net40 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net47 cn net87 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net40 net47 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net48 c net47 VNW PHVT11LL_CKT W=0.37u L=40.00n
XX1 net48 D VDD VNW PHVT11LL_CKT W=0.47u L=40.00n
.ENDS DQV8_12TH40
.SUBCKT DRNQNV0_12TH40 CK D QN RDN VDD VSS
XX21 net147 net152 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net152 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX29 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX26 net88 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX24 net112 R VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX1 net177 D VDD VNW PHVT11LL_CKT W=0.21u L=40.00n
XX0 net177 c net0152 VNW PHVT11LL_CKT W=0.21u L=40.00n
XX5 net169 net0152 net112 VNW PHVT11LL_CKT W=0.44u L=40.00n
XX7 net0152 cn net108 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net108 net169 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.38u L=40.00n
XX15 net169 cn net152 VNW PHVT11LL_CKT W=0.28u L=40.00n
XX19 net84 net147 net88 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net152 c net84 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX25 net169 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX28 R RDN VSS VPW NHVT11LL_CKT W=210.00n L=40.00n
XX27 net152 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net177 D VSS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX3 net177 cn net0152 VPW NHVT11LL_CKT W=0.28u L=40.00n
XX4 net169 net0152 VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX6 net0152 c net161 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net161 net169 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX14 net169 c net152 VPW NHVT11LL_CKT W=0.26u L=40.00n
XX16 net145 net147 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net152 cn net145 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net147 net152 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net152 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
.ENDS DRNQNV0_12TH40
.SUBCKT DRNQNV2_12TH40 CK D QN RDN VDD VSS
XX25 net84 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX28 R RDN VSS VPW NHVT11LL_CKT W=210.00n L=40.00n
XX27 net99 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net100 D VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX3 net100 cn net092 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX4 net84 net092 VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX6 net092 c net92 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net92 net84 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=190.00n L=40.00n
XX14 net84 c net99 VPW NHVT11LL_CKT W=0.28u L=40.00n
XX16 net72 net74 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net99 cn net72 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net74 net99 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net99 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX29 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX26 net19 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX24 net31 R VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX1 net100 D VDD VNW PHVT11LL_CKT W=0.27u L=40.00n
XX0 net100 c net092 VNW PHVT11LL_CKT W=0.27u L=40.00n
XX5 net84 net092 net31 VNW PHVT11LL_CKT W=0.55u L=40.00n
XX7 net092 cn net35 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net35 net84 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX15 net84 cn net99 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX19 net23 net74 net19 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net99 c net23 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net74 net99 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net99 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS DRNQNV2_12TH40
.SUBCKT DRNQNV4_12TH40 CK D QN RDN VDD VSS
XX21 net147 net152 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net152 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX29 R RDN VDD VNW PHVT11LL_CKT W=0.3u L=40.00n
XX26 net88 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX24 net112 R VDD VNW PHVT11LL_CKT W=0.91u L=40.00n
XX1 net177 D VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX0 net177 c net0152 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX5 net169 net0152 net112 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX7 net0152 cn net108 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net108 net169 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX15 net169 cn net152 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX19 net84 net147 net88 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net152 c net84 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX25 net169 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX28 R RDN VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX27 net152 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net177 D VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX3 net177 cn net0152 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX4 net169 net0152 VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX6 net0152 c net161 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net161 net169 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=190.00n L=40.00n
XX14 net169 c net152 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX16 net145 net147 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net152 cn net145 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net147 net152 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net152 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
.ENDS DRNQNV4_12TH40
.SUBCKT DRNQNV6_12TH40 CK D QN RDN VDD VSS
XX21 net147 net152 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net152 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX29 R RDN VDD VNW PHVT11LL_CKT W=0.3u L=40.00n
XX26 net88 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX24 net112 R VDD VNW PHVT11LL_CKT W=0.91u L=40.00n
XX1 net177 D VDD VNW PHVT11LL_CKT W=0.37u L=40.00n
XX0 net177 c net0152 VNW PHVT11LL_CKT W=0.37u L=40.00n
XX5 net169 net0152 net112 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX7 net0152 cn net108 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net108 net169 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.21u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.3u L=40.00n
XX15 net169 cn net152 VNW PHVT11LL_CKT W=0.49u L=40.00n
XX19 net84 net147 net88 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net152 c net84 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX25 net169 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX28 R RDN VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX27 net152 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net177 D VSS VPW NHVT11LL_CKT W=0.59u L=40.00n
XX3 net177 cn net0152 VPW NHVT11LL_CKT W=0.5u L=40.00n
XX4 net169 net0152 VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX6 net0152 c net161 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net161 net169 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX14 net169 c net152 VPW NHVT11LL_CKT W=0.27u L=40.00n
XX16 net145 net147 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net152 cn net145 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net147 net152 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net152 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
.ENDS DRNQNV6_12TH40
.SUBCKT DRNQV0_12TH40 CK D Q RDN VDD VSS
XX28 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX26 net52 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX24 net28 R VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX1 net77 D VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX0 net77 c net0151 VNW PHVT11LL_CKT W=0.22u L=40.00n
XX5 net85 net0151 net28 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX7 net0151 cn net32 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net32 net85 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX15 net85 cn net108 VNW PHVT11LL_CKT W=0.23u L=40.00n
XX19 net56 net111 net52 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net108 c net56 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net111 net108 VDD VNW PHVT11LL_CKT W=0.21u L=40.00n
XX23 Q net111 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX29 R RDN VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX25 net85 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX27 net108 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net77 D VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX3 net77 cn net0151 VPW NHVT11LL_CKT W=0.31u L=40.00n
XX4 net85 net0151 VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX6 net0151 c net93 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net93 net85 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX14 net85 c net108 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX16 net109 net111 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net108 cn net109 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net111 net108 VSS VPW NHVT11LL_CKT W=0.195u L=40.00n
XX22 Q net111 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
.ENDS DRNQV0_12TH40
.SUBCKT DRNQV2_12TH40 CK D Q RDN VDD VSS
XX28 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX26 net52 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX24 net28 R VDD VNW PHVT11LL_CKT W=460.00n L=40.00n
XX1 net77 D VDD VNW PHVT11LL_CKT W=0.24u L=40.00n
XX0 net77 c net0151 VNW PHVT11LL_CKT W=0.24u L=40.00n
XX5 net85 net0151 net28 VNW PHVT11LL_CKT W=460.00n L=40.00n
XX7 net0151 cn net32 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net32 net85 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX15 net85 cn net108 VNW PHVT11LL_CKT W=0.29u L=40.00n
XX19 net56 net111 net52 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net108 c net56 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net111 net108 VDD VNW PHVT11LL_CKT W=0.345u L=40.00n
XX23 Q net111 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX29 R RDN VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX25 net85 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX27 net108 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net77 D VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX3 net77 cn net0151 VPW NHVT11LL_CKT W=0.31u L=40.00n
XX4 net85 net0151 VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX6 net0151 c net93 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net93 net85 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX14 net85 c net108 VPW NHVT11LL_CKT W=0.28u L=40.00n
XX16 net109 net111 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net108 cn net109 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net111 net108 VSS VPW NHVT11LL_CKT W=325.00n L=40.00n
XX22 Q net111 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
.ENDS DRNQV2_12TH40
.SUBCKT DRNQV4_12TH40 CK D Q RDN VDD VSS
XX28 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX26 net52 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX24 net28 R VDD VNW PHVT11LL_CKT W=0.91u L=40.00n
XX1 net77 D VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX0 net77 c net0151 VNW PHVT11LL_CKT W=0.31u L=40.00n
XX5 net85 net0151 net28 VNW PHVT11LL_CKT W=0.52u L=40.00n
XX7 net0151 cn net32 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net32 net85 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX15 net85 cn net108 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX19 net56 net111 net52 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net108 c net56 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net111 net108 VDD VNW PHVT11LL_CKT W=0.535u L=40.00n
XX23 Q net111 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX29 R RDN VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX25 net85 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX27 net108 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net77 D VSS VPW NHVT11LL_CKT W=0.46u L=40.00n
XX3 net77 cn net0151 VPW NHVT11LL_CKT W=0.37u L=40.00n
XX4 net85 net0151 VSS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX6 net0151 c net93 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net93 net85 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX14 net85 c net108 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX16 net109 net111 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net108 cn net109 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net111 net108 VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX22 Q net111 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
.ENDS DRNQV4_12TH40
.SUBCKT DRNQV6_12TH40 CK D Q RDN VDD VSS
XX28 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX26 net52 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX24 net28 R VDD VNW PHVT11LL_CKT W=0.81u L=40.00n
XX1 net77 D VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX0 net77 c net0151 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX5 net85 net0151 net28 VNW PHVT11LL_CKT W=0.56u L=40.00n
XX7 net0151 cn net32 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net32 net85 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
XX15 net85 cn net108 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX19 net56 net111 net52 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net108 c net56 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net111 net108 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX23 Q net111 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX29 R RDN VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX25 net85 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX27 net108 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net77 D VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX3 net77 cn net0151 VPW NHVT11LL_CKT W=0.42u L=40.00n
XX4 net85 net0151 VSS VPW NHVT11LL_CKT W=0.44u L=40.00n
XX6 net0151 c net93 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net93 net85 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX14 net85 c net108 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX16 net109 net111 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net108 cn net109 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net111 net108 VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX22 Q net111 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
.ENDS DRNQV6_12TH40
.SUBCKT DRNQV8_12TH40 CK D Q RDN VDD VSS
XX28 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX26 net52 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX24 net28 R VDD VNW PHVT11LL_CKT W=0.91u L=40.00n
XX1 net77 D VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX0 net77 c net0151 VNW PHVT11LL_CKT W=0.35u L=40.00n
XX5 net85 net0151 net28 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX7 net0151 cn net32 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net32 net85 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.21u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
XX15 net85 cn net108 VNW PHVT11LL_CKT W=0.49u L=40.00n
XX19 net56 net111 net52 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net108 c net56 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net111 net108 VDD VNW PHVT11LL_CKT W=0.68u L=40.00n
XX23 Q net111 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX29 R RDN VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX25 net85 R VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX27 net108 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net77 D VSS VPW NHVT11LL_CKT W=0.59u L=40.00n
XX3 net77 cn net0151 VPW NHVT11LL_CKT W=0.5u L=40.00n
XX4 net85 net0151 VSS VPW NHVT11LL_CKT W=0.42u L=40.00n
XX6 net0151 c net93 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net93 net85 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX14 net85 c net108 VPW NHVT11LL_CKT W=0.42u L=40.00n
XX16 net109 net111 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net108 cn net109 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net111 net108 VSS VPW NHVT11LL_CKT W=0.72u L=40.00n
XX22 Q net111 VSS VPW NHVT11LL_CKT W=2.14u L=40.00n
.ENDS DRNQV8_12TH40
.SUBCKT DRSNQNV0_12TH40 CK D QN RDN SDN VDD VSS
XX33 R RDN VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX22 QN net23 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX18 net18 net23 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net23 cn net16 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX16 net16 net18 net60 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX14 net40 c net23 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX9 net32 net40 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net47 c net32 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net40 net47 net52 VPW NHVT11LL_CKT W=0.26u L=40.00n
XX3 net48 cn net47 VPW NHVT11LL_CKT W=0.28u L=40.00n
XX2 net48 D VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX26 net52 SDN VSS VPW NHVT11LL_CKT W=0.36u L=40.00n
XX27 net40 R net52 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX29 net60 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX31 net23 SDN net68 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX32 net68 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX34 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX23 QN net23 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX21 net18 net23 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net23 c net83 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX19 net83 net18 net87 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX15 net40 cn net23 VNW PHVT11LL_CKT W=0.285u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX8 net107 net40 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net47 cn net107 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net40 net47 net111 VNW PHVT11LL_CKT W=0.39u L=40.00n
XX0 net48 c net47 VNW PHVT11LL_CKT W=0.22u L=40.00n
XX1 net48 D VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX24 net40 SDN VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX25 net111 R VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
XX28 net87 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX30 net23 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS DRSNQNV0_12TH40
.SUBCKT DRSNQNV2_12TH40 CK D QN RDN SDN VDD VSS
XX33 R RDN VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX22 QN net23 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX18 net18 net23 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net23 cn net16 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX16 net16 net18 net60 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX14 net40 c net23 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX9 net32 net40 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net47 c net32 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net40 net47 net52 VPW NHVT11LL_CKT W=0.27u L=40.00n
XX3 net48 cn net47 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX2 net48 D VSS VPW NHVT11LL_CKT W=0.355u L=40.00n
XX26 net52 SDN VSS VPW NHVT11LL_CKT W=0.46u L=40.00n
XX27 net40 R net52 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX29 net60 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX31 net23 SDN net68 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX32 net68 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX34 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX23 QN net23 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX21 net18 net23 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net23 c net83 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX19 net83 net18 net87 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX15 net40 cn net23 VNW PHVT11LL_CKT W=0.31u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX8 net107 net40 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net47 cn net107 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net40 net47 net111 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX0 net48 c net47 VNW PHVT11LL_CKT W=0.28u L=40.00n
XX1 net48 D VDD VNW PHVT11LL_CKT W=0.28u L=40.00n
XX24 net40 SDN VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX25 net111 R VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX28 net87 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX30 net23 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS DRSNQNV2_12TH40
.SUBCKT DRSNQNV4_12TH40 CK D QN RDN SDN VDD VSS
XX33 R RDN VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX22 QN net23 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX18 net18 net23 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net23 cn net16 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX16 net16 net18 net60 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX14 net40 c net23 VPW NHVT11LL_CKT W=0.29u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX9 net32 net40 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net47 c net32 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net40 net47 net52 VPW NHVT11LL_CKT W=0.32u L=40.00n
XX3 net48 cn net47 VPW NHVT11LL_CKT W=0.34u L=40.00n
XX2 net48 D VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX26 net52 SDN VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX27 net40 R net52 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX29 net60 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX31 net23 SDN net68 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX32 net68 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX34 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX23 QN net23 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX21 net18 net23 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net23 c net83 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX19 net83 net18 net87 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX15 net40 cn net23 VNW PHVT11LL_CKT W=0.425u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX8 net107 net40 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net47 cn net107 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net40 net47 net111 VNW PHVT11LL_CKT W=0.545u L=40.00n
XX0 net48 c net47 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX1 net48 D VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX24 net40 SDN VDD VNW PHVT11LL_CKT W=0.21u L=40.00n
XX25 net111 R VDD VNW PHVT11LL_CKT W=0.78u L=40.00n
XX28 net87 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX30 net23 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS DRSNQNV4_12TH40
.SUBCKT DRSNQNV6_12TH40 CK D QN RDN SDN VDD VSS
XX33 R RDN VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX22 QN net23 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX18 net18 net23 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net23 cn net16 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX16 net16 net18 net60 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX14 net40 c net23 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX9 net32 net40 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net47 c net32 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net40 net47 net52 VPW NHVT11LL_CKT W=0.34u L=40.00n
XX3 net48 cn net47 VPW NHVT11LL_CKT W=0.42u L=40.00n
XX2 net48 D VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX26 net52 SDN VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX27 net40 R net52 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX29 net60 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX31 net23 SDN net68 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX32 net68 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX34 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX23 QN net23 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX21 net18 net23 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net23 c net83 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX19 net83 net18 net87 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX15 net40 cn net23 VNW PHVT11LL_CKT W=0.49u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX8 net107 net40 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net47 cn net107 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net40 net47 net111 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net48 c net47 VNW PHVT11LL_CKT W=0.42u L=40.00n
XX1 net48 D VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX24 net40 SDN VDD VNW PHVT11LL_CKT W=0.21u L=40.00n
XX25 net111 R VDD VNW PHVT11LL_CKT W=0.91u L=40.00n
XX28 net87 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX30 net23 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS DRSNQNV6_12TH40
.SUBCKT DRSNQV0_12TH40 CK D Q RDN SDN VDD VSS
XX33 R RDN VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX22 Q net18 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX18 net18 net23 VSS VPW NHVT11LL_CKT W=0.195u L=40.00n
XX17 net23 cn net16 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX16 net16 net18 net60 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX14 net40 c net23 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX9 net32 net40 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net47 c net32 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net40 net47 net52 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX3 net48 cn net47 VPW NHVT11LL_CKT W=0.28u L=40.00n
XX2 net48 D VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX26 net52 SDN VSS VPW NHVT11LL_CKT W=0.36u L=40.00n
XX27 net40 R net52 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX29 net60 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX31 net23 SDN net68 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX32 net68 R VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX34 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX23 Q net18 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX21 net18 net23 VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX20 net23 c net83 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX19 net83 net18 net87 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX15 net40 cn net23 VNW PHVT11LL_CKT W=0.255u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.38u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX8 net107 net40 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net47 cn net107 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net40 net47 net111 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX0 net48 c net47 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX1 net48 D VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX24 net40 SDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX25 net111 R VDD VNW PHVT11LL_CKT W=470.00n L=40.00n
XX28 net87 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX30 net23 SDN VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
.ENDS DRSNQV0_12TH40
.SUBCKT DRSNQV2_12TH40 CK D Q RDN SDN VDD VSS
XX33 R RDN VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX22 Q net18 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX18 net18 net23 VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX17 net23 cn net16 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX16 net16 net18 net60 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX14 net40 c net23 VPW NHVT11LL_CKT W=0.27u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX9 net32 net40 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net47 c net32 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net40 net47 net52 VPW NHVT11LL_CKT W=390.00n L=40.00n
XX3 net48 cn net47 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX2 net48 D VSS VPW NHVT11LL_CKT W=0.39u L=40.00n
XX26 net52 SDN VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX27 net40 R net52 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX29 net60 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX31 net23 SDN net68 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX32 net68 R VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX34 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX23 Q net18 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX21 net18 net23 VDD VNW PHVT11LL_CKT W=350.00n L=40.00n
XX20 net23 c net83 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX19 net83 net18 net87 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX15 net40 cn net23 VNW PHVT11LL_CKT W=0.41u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.38u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX8 net107 net40 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net47 cn net107 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net40 net47 net111 VNW PHVT11LL_CKT W=0.51u L=40.00n
XX0 net48 c net47 VNW PHVT11LL_CKT W=0.27u L=40.00n
XX1 net48 D VDD VNW PHVT11LL_CKT W=0.27u L=40.00n
XX24 net40 SDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX25 net111 R VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX28 net87 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX30 net23 SDN VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
.ENDS DRSNQV2_12TH40
.SUBCKT DRSNQV4_12TH40 CK D Q RDN SDN VDD VSS
XX33 R RDN VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX22 Q net18 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX18 net18 net23 VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX17 net23 cn net16 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX16 net16 net18 net60 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX14 net40 c net23 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX9 net32 net40 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net47 c net32 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net40 net47 net52 VPW NHVT11LL_CKT W=0.45u L=40.00n
XX3 net48 cn net47 VPW NHVT11LL_CKT W=0.34u L=40.00n
XX2 net48 D VSS VPW NHVT11LL_CKT W=0.395u L=40.00n
XX26 net52 SDN VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX27 net40 R net52 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX29 net60 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX31 net23 SDN net68 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX32 net68 R VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX34 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX23 Q net18 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX21 net18 net23 VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX20 net23 c net83 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX19 net83 net18 net87 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX15 net40 cn net23 VNW PHVT11LL_CKT W=0.385u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX8 net107 net40 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net47 cn net107 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net40 net47 net111 VNW PHVT11LL_CKT W=0.505u L=40.00n
XX0 net48 c net47 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX1 net48 D VDD VNW PHVT11LL_CKT W=0.3u L=40.00n
XX24 net40 SDN VDD VNW PHVT11LL_CKT W=0.21u L=40.00n
XX25 net111 R VDD VNW PHVT11LL_CKT W=0.91u L=40.00n
XX28 net87 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX30 net23 SDN VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
.ENDS DRSNQV4_12TH40
.SUBCKT DRSNQV6_12TH40 CK D Q RDN SDN VDD VSS
XX33 R RDN VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX22 Q net18 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX18 net18 net23 VSS VPW NHVT11LL_CKT W=0.51u L=40.00n
XX17 net23 cn net16 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX16 net16 net18 net60 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX14 net40 c net23 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX9 net32 net40 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net47 c net32 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net40 net47 net52 VPW NHVT11LL_CKT W=0.5u L=40.00n
XX3 net48 cn net47 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX2 net48 D VSS VPW NHVT11LL_CKT W=0.52u L=40.00n
XX26 net52 SDN VSS VPW NHVT11LL_CKT W=0.48u L=40.00n
XX27 net40 R net52 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX29 net60 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX31 net23 SDN net68 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX32 net68 R VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX34 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX23 Q net18 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX21 net18 net23 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX20 net23 c net83 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX19 net83 net18 net87 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX15 net40 cn net23 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX8 net107 net40 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net47 cn net107 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net40 net47 net111 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net48 c net47 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX1 net48 D VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX24 net40 SDN VDD VNW PHVT11LL_CKT W=0.21u L=40.00n
XX25 net111 R VDD VNW PHVT11LL_CKT W=0.91u L=40.00n
XX28 net87 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX30 net23 SDN VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
.ENDS DRSNQV6_12TH40
.SUBCKT DRSNQV8_12TH40 CK D Q RDN SDN VDD VSS
XX33 R RDN VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX22 Q net18 VSS VPW NHVT11LL_CKT W=2.14u L=40.00n
XX18 net18 net23 VSS VPW NHVT11LL_CKT W=0.68u L=40.00n
XX17 net23 cn net16 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX16 net16 net18 net60 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX14 net40 c net23 VPW NHVT11LL_CKT W=0.48u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX9 net32 net40 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net47 c net32 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net40 net47 net52 VPW NHVT11LL_CKT W=0.48u L=40.00n
XX3 net48 cn net47 VPW NHVT11LL_CKT W=0.5u L=40.00n
XX2 net48 D VSS VPW NHVT11LL_CKT W=0.59u L=40.00n
XX26 net52 SDN VSS VPW NHVT11LL_CKT W=0.48u L=40.00n
XX27 net40 R net52 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX29 net60 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX31 net23 SDN net68 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX32 net68 R VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX34 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX23 Q net18 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX21 net18 net23 VDD VNW PHVT11LL_CKT W=0.7u L=40.00n
XX20 net23 c net83 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX19 net83 net18 net87 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX15 net40 cn net23 VNW PHVT11LL_CKT W=0.52u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX8 net107 net40 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net47 cn net107 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net40 net47 net111 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net48 c net47 VNW PHVT11LL_CKT W=0.44u L=40.00n
XX1 net48 D VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX24 net40 SDN VDD VNW PHVT11LL_CKT W=0.21u L=40.00n
XX25 net111 R VDD VNW PHVT11LL_CKT W=0.91u L=40.00n
XX28 net87 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX30 net23 SDN VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
.ENDS DRSNQV8_12TH40
.SUBCKT DSNQNV0_12TH40 CK D QN SDN VDD VSS
XX24 net36 SDN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX22 QN net27 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX18 net14 net27 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net27 cn net12 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX16 net12 net14 net4 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX14 net48 c net27 VPW NHVT11LL_CKT W=0.24u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net28 net48 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net55 c net28 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net48 net55 net36 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX3 net56 cn net55 VPW NHVT11LL_CKT W=0.22u L=40.00n
XX2 net56 D VSS VPW NHVT11LL_CKT W=0.36u L=40.00n
XX25 net4 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX28 net48 SDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX29 net27 SDN VDD VNW PHVT11LL_CKT W=0.16u L=40.00n
XX23 QN net27 VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX21 net14 net27 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net27 c net63 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net63 net14 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net48 cn net27 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net91 net48 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net55 cn net91 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net48 net55 VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX0 net56 c net55 VNW PHVT11LL_CKT W=0.22u L=40.00n
XX1 net56 D VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
.ENDS DSNQNV0_12TH40
.SUBCKT DSNQNV2_12TH40 CK D QN SDN VDD VSS
XX24 net36 SDN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX22 QN net27 VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX18 net14 net27 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net27 cn net12 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX16 net12 net14 net4 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX14 net48 c net27 VPW NHVT11LL_CKT W=330.00n L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=190.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX9 net28 net48 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net55 c net28 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net48 net55 net36 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX3 net56 cn net55 VPW NHVT11LL_CKT W=330.00n L=40.00n
XX2 net56 D VSS VPW NHVT11LL_CKT W=0.44u L=40.00n
XX25 net4 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX28 net48 SDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX29 net27 SDN VDD VNW PHVT11LL_CKT W=0.16u L=40.00n
XX23 QN net27 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX21 net14 net27 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net27 c net63 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net63 net14 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net48 cn net27 VNW PHVT11LL_CKT W=0.29u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.13u L=40.00n
XX8 net91 net48 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net55 cn net91 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net48 net55 VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX0 net56 c net55 VNW PHVT11LL_CKT W=0.25u L=40.00n
XX1 net56 D VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
.ENDS DSNQNV2_12TH40
.SUBCKT DSNQNV4_12TH40 CK D QN SDN VDD VSS
XX24 net36 SDN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX22 QN net27 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX18 net14 net27 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net27 cn net12 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX16 net12 net14 net4 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX14 net48 c net27 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX9 net28 net48 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net55 c net28 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net48 net55 net36 VPW NHVT11LL_CKT W=0.61u L=40.00n
XX3 net56 cn net55 VPW NHVT11LL_CKT W=0.435u L=40.00n
XX2 net56 D VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX25 net4 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX28 net48 SDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX29 net27 SDN VDD VNW PHVT11LL_CKT W=0.16u L=40.00n
XX23 QN net27 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX21 net14 net27 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net27 c net63 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net63 net14 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net48 cn net27 VNW PHVT11LL_CKT W=0.4u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX8 net91 net48 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net55 cn net91 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net48 net55 VDD VNW PHVT11LL_CKT W=0.49u L=40.00n
XX0 net56 c net55 VNW PHVT11LL_CKT W=0.32u L=40.00n
XX1 net56 D VDD VNW PHVT11LL_CKT W=0.32u L=40.00n
.ENDS DSNQNV4_12TH40
.SUBCKT DSNQNV6_12TH40 CK D QN SDN VDD VSS
XX24 net36 SDN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX22 QN net27 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX18 net14 net27 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net27 cn net12 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX16 net12 net14 net4 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX14 net48 c net27 VPW NHVT11LL_CKT W=0.48u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX9 net28 net48 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net55 c net28 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net48 net55 net36 VPW NHVT11LL_CKT W=0.61u L=40.00n
XX3 net56 cn net55 VPW NHVT11LL_CKT W=0.45u L=40.00n
XX2 net56 D VSS VPW NHVT11LL_CKT W=0.59u L=40.00n
XX25 net4 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX28 net48 SDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX29 net27 SDN VDD VNW PHVT11LL_CKT W=0.16u L=40.00n
XX23 QN net27 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX21 net14 net27 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net27 c net63 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net63 net14 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net48 cn net27 VNW PHVT11LL_CKT W=0.49u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.21u L=40.00n
XX8 net91 net48 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net55 cn net91 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net48 net55 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net56 c net55 VNW PHVT11LL_CKT W=0.42u L=40.00n
XX1 net56 D VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
.ENDS DSNQNV6_12TH40
.SUBCKT DSNQV0_12TH40 CK D Q SDN VDD VSS
XX2 net64 D VSS VPW NHVT11LL_CKT W=0.425u L=40.00n
XX3 net64 cn net71 VPW NHVT11LL_CKT W=0.22u L=40.00n
XX4 net72 net71 net84 VPW NHVT11LL_CKT W=0.32u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX24 net84 SDN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX6 net71 c net92 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net92 net72 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net72 c net99 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX18 net106 net99 VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX22 Q net106 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX16 net104 net106 net112 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net99 cn net104 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX25 net112 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX1 net64 D VDD VNW PHVT11LL_CKT W=0.26u L=40.00n
XX0 net64 c net71 VNW PHVT11LL_CKT W=260.00n L=40.00n
XX5 net72 net71 VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.38u L=40.00n
XX28 net72 SDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX7 net71 cn net35 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net35 net72 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net72 cn net99 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX21 net106 net99 VDD VNW PHVT11LL_CKT W=0.27u L=40.00n
XX23 Q net106 VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX29 net99 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net59 net106 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net99 c net59 VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS DSNQV0_12TH40
.SUBCKT DSNQV2_12TH40 CK D Q SDN VDD VSS
XX2 net64 D VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX3 net64 cn net71 VPW NHVT11LL_CKT W=0.295u L=40.00n
XX4 net72 net71 net84 VPW NHVT11LL_CKT W=0.45u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=130.00n L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=185.00n L=40.00n
XX24 net84 SDN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX6 net71 c net92 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net92 net72 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net72 c net99 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX18 net106 net99 VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX22 Q net106 VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX16 net104 net106 net112 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net99 cn net104 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX25 net112 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX1 net64 D VDD VNW PHVT11LL_CKT W=0.26u L=40.00n
XX0 net64 c net71 VNW PHVT11LL_CKT W=260.00n L=40.00n
XX5 net72 net71 VDD VNW PHVT11LL_CKT W=0.47u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX28 net72 SDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX7 net71 cn net35 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net35 net72 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net72 cn net99 VNW PHVT11LL_CKT W=0.295u L=40.00n
XX21 net106 net99 VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX23 Q net106 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX29 net99 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net59 net106 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net99 c net59 VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS DSNQV2_12TH40
.SUBCKT DSNQV4_12TH40 CK D Q SDN VDD VSS
XX2 net64 D VSS VPW NHVT11LL_CKT W=0.48u L=40.00n
XX3 net64 cn net71 VPW NHVT11LL_CKT W=0.35u L=40.00n
XX4 net72 net71 net84 VPW NHVT11LL_CKT W=0.475u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX24 net84 SDN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX6 net71 c net92 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net92 net72 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net72 c net99 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX18 net106 net99 VSS VPW NHVT11LL_CKT W=0.325u L=40.00n
XX22 Q net106 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX16 net104 net106 net112 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net99 cn net104 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX25 net112 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX1 net64 D VDD VNW PHVT11LL_CKT W=0.32u L=40.00n
XX0 net64 c net71 VNW PHVT11LL_CKT W=0.28u L=40.00n
XX5 net72 net71 VDD VNW PHVT11LL_CKT W=0.48u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.18u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX28 net72 SDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX7 net71 cn net35 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net35 net72 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net72 cn net99 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX21 net106 net99 VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX23 Q net106 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX29 net99 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net59 net106 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net99 c net59 VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS DSNQV4_12TH40
.SUBCKT DSNQV6_12TH40 CK D Q SDN VDD VSS
XX2 net64 D VSS VPW NHVT11LL_CKT W=0.57u L=40.00n
XX3 net64 cn net71 VPW NHVT11LL_CKT W=0.42u L=40.00n
XX4 net72 net71 net84 VPW NHVT11LL_CKT W=0.61u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX24 net84 SDN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX6 net71 c net92 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net92 net72 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net72 c net99 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX18 net106 net99 VSS VPW NHVT11LL_CKT W=0.42u L=40.00n
XX22 Q net106 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX16 net104 net106 net112 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net99 cn net104 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX25 net112 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX1 net64 D VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX0 net64 c net71 VNW PHVT11LL_CKT W=0.32u L=40.00n
XX5 net72 net71 VDD VNW PHVT11LL_CKT W=0.55u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX28 net72 SDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX7 net71 cn net35 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net35 net72 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net72 cn net99 VNW PHVT11LL_CKT W=0.37u L=40.00n
XX21 net106 net99 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX23 Q net106 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX29 net99 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net59 net106 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net99 c net59 VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS DSNQV6_12TH40
.SUBCKT DSNQV8_12TH40 CK D Q SDN VDD VSS
XX2 net64 D VSS VPW NHVT11LL_CKT W=0.59u L=40.00n
XX3 net64 cn net71 VPW NHVT11LL_CKT W=0.5u L=40.00n
XX4 net72 net71 net84 VPW NHVT11LL_CKT W=0.61u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX24 net84 SDN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX6 net71 c net92 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net92 net72 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net72 c net99 VPW NHVT11LL_CKT W=0.49u L=40.00n
XX18 net106 net99 VSS VPW NHVT11LL_CKT W=0.63u L=40.00n
XX22 Q net106 VSS VPW NHVT11LL_CKT W=2.14u L=40.00n
XX16 net104 net106 net112 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net99 cn net104 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX25 net112 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX1 net64 D VDD VNW PHVT11LL_CKT W=0.47u L=40.00n
XX0 net64 c net71 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX5 net72 net71 VDD VNW PHVT11LL_CKT W=0.53u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.21u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX28 net72 SDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX7 net71 cn net35 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net35 net72 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net72 cn net99 VNW PHVT11LL_CKT W=0.49u L=40.00n
XX21 net106 net99 VDD VNW PHVT11LL_CKT W=0.93u L=40.00n
XX23 Q net106 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX29 net99 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net59 net106 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net99 c net59 VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS DSNQV8_12TH40
.SUBCKT DXQNV2_12TH40 CK DA DB QN SA VDD VSS
XX43 net140 SAN net171 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX6 net103 c net108 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX3 net156 cn net103 VPW NHVT11LL_CKT W=0.29u L=40.00n
XX4 net104 net103 VSS VPW NHVT11LL_CKT W=355.00n L=40.00n
XX9 net108 net104 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=130.00n L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=185.00n L=40.00n
XX14 net104 c net123 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX16 net124 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net123 cn net124 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 s net123 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX22 QN s VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX26 net140 DB VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX24 SAN SA VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX34 net156 net171 VSS VPW NHVT11LL_CKT W=0.435u L=40.00n
XX45 net172 SA net171 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX46 net172 DA VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX0 net156 c net103 VNW PHVT11LL_CKT W=0.24u L=40.00n
XX5 net104 net103 VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX7 net103 cn net19 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net19 net104 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX15 net104 cn net123 VNW PHVT11LL_CKT W=260.00n L=40.00n
XX19 net43 s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net123 c net43 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX21 s net123 VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX23 QN s VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX44 net140 SA net171 VNW PHVT11LL_CKT W=0.35u L=40.00n
XX25 SAN SA VDD VNW PHVT11LL_CKT W=315.00n L=40.00n
XX27 net140 DB VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX35 net156 net171 VDD VNW PHVT11LL_CKT W=0.24u L=40.00n
XX47 net172 SAN net171 VNW PHVT11LL_CKT W=0.35u L=40.00n
XX48 net172 DA VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
.ENDS DXQNV2_12TH40
.SUBCKT DXQNV4_12TH40 CK DA DB QN SA VDD VSS
XX43 net140 SAN net171 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX6 net103 c net108 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX3 net156 cn net103 VPW NHVT11LL_CKT W=0.29u L=40.00n
XX4 net104 net103 VSS VPW NHVT11LL_CKT W=0.385u L=40.00n
XX9 net108 net104 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=130.00n L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=185.00n L=40.00n
XX14 net104 c net123 VPW NHVT11LL_CKT W=0.29u L=40.00n
XX16 net124 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net123 cn net124 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 s net123 VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX22 QN s VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX26 net140 DB VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX24 SAN SA VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX34 net156 net171 VSS VPW NHVT11LL_CKT W=0.495u L=40.00n
XX45 net172 SA net171 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX46 net172 DA VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX0 net156 c net103 VNW PHVT11LL_CKT W=0.24u L=40.00n
XX5 net104 net103 VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX7 net103 cn net19 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net19 net104 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX15 net104 cn net123 VNW PHVT11LL_CKT W=260.00n L=40.00n
XX19 net43 s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net123 c net43 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX21 s net123 VDD VNW PHVT11LL_CKT W=0.51u L=40.00n
XX23 QN s VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX44 net140 SA net171 VNW PHVT11LL_CKT W=0.35u L=40.00n
XX25 SAN SA VDD VNW PHVT11LL_CKT W=315.00n L=40.00n
XX27 net140 DB VDD VNW PHVT11LL_CKT W=0.55u L=40.00n
XX35 net156 net171 VDD VNW PHVT11LL_CKT W=0.24u L=40.00n
XX47 net172 SAN net171 VNW PHVT11LL_CKT W=0.35u L=40.00n
XX48 net172 DA VDD VNW PHVT11LL_CKT W=0.55u L=40.00n
.ENDS DXQNV4_12TH40
.SUBCKT DXQNV6_12TH40 CK DA DB QN SA VDD VSS
XX43 net140 SAN net171 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX6 net103 c net108 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX3 net156 cn net103 VPW NHVT11LL_CKT W=0.29u L=40.00n
XX4 net104 net103 VSS VPW NHVT11LL_CKT W=0.385u L=40.00n
XX9 net108 net104 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=130.00n L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=185.00n L=40.00n
XX14 net104 c net123 VPW NHVT11LL_CKT W=0.29u L=40.00n
XX16 net124 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net123 cn net124 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 s net123 VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX22 QN s VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX26 net140 DB VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX24 SAN SA VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX34 net156 net171 VSS VPW NHVT11LL_CKT W=0.495u L=40.00n
XX45 net172 SA net171 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX46 net172 DA VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX0 net156 c net103 VNW PHVT11LL_CKT W=0.24u L=40.00n
XX5 net104 net103 VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX7 net103 cn net19 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net19 net104 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX15 net104 cn net123 VNW PHVT11LL_CKT W=260.00n L=40.00n
XX19 net43 s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net123 c net43 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX21 s net123 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX23 QN s VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX44 net140 SA net171 VNW PHVT11LL_CKT W=0.35u L=40.00n
XX25 SAN SA VDD VNW PHVT11LL_CKT W=315.00n L=40.00n
XX27 net140 DB VDD VNW PHVT11LL_CKT W=0.55u L=40.00n
XX35 net156 net171 VDD VNW PHVT11LL_CKT W=0.24u L=40.00n
XX47 net172 SAN net171 VNW PHVT11LL_CKT W=0.35u L=40.00n
XX48 net172 DA VDD VNW PHVT11LL_CKT W=0.55u L=40.00n
.ENDS DXQNV6_12TH40
.SUBCKT DXQV2_12TH40 CK DA DB Q SA VDD VSS
XX43 net140 SAN net171 VPW NHVT11LL_CKT W=0.19u L=40.00n
XX6 net103 c net108 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX3 net156 cn net103 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX4 net104 net103 VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX9 net108 net104 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX14 net104 c net123 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX16 net124 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net123 cn net124 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 s net123 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX22 Q net123 VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX26 net140 DB VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX24 SAN SA VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX34 net156 net171 VSS VPW NHVT11LL_CKT W=0.49u L=40.00n
XX45 net172 SA net171 VPW NHVT11LL_CKT W=0.19u L=40.00n
XX46 net172 DA VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX0 net156 c net103 VNW PHVT11LL_CKT W=0.25u L=40.00n
XX5 net104 net103 VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX7 net103 cn net19 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net19 net104 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX15 net104 cn net123 VNW PHVT11LL_CKT W=0.27u L=40.00n
XX19 net43 s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net123 c net43 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX21 s net123 VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX23 Q net123 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX44 net140 SA net171 VNW PHVT11LL_CKT W=0.405u L=40.00n
XX25 SAN SA VDD VNW PHVT11LL_CKT W=0.34u L=40.00n
XX27 net140 DB VDD VNW PHVT11LL_CKT W=0.55u L=40.00n
XX35 net156 net171 VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX47 net172 SAN net171 VNW PHVT11LL_CKT W=0.405u L=40.00n
XX48 net172 DA VDD VNW PHVT11LL_CKT W=0.55u L=40.00n
.ENDS DXQV2_12TH40
.SUBCKT DXQV4_12TH40 CK DA DB Q SA VDD VSS
XX43 net140 SAN net171 VPW NHVT11LL_CKT W=0.21u L=40.00n
XX6 net103 c net108 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX3 net156 cn net103 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX4 net104 net103 VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX9 net108 net104 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=130.00n L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX14 net104 c net123 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX16 net124 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net123 cn net124 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 s net123 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX22 Q net123 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX26 net140 DB VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX24 SAN SA VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX34 net156 net171 VSS VPW NHVT11LL_CKT W=0.49u L=40.00n
XX45 net172 SA net171 VPW NHVT11LL_CKT W=0.21u L=40.00n
XX46 net172 DA VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX0 net156 c net103 VNW PHVT11LL_CKT W=0.25u L=40.00n
XX5 net104 net103 VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX7 net103 cn net19 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net19 net104 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX15 net104 cn net123 VNW PHVT11LL_CKT W=0.37u L=40.00n
XX19 net43 s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net123 c net43 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX21 s net123 VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX23 Q net123 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX44 net140 SA net171 VNW PHVT11LL_CKT W=0.455u L=40.00n
XX25 SAN SA VDD VNW PHVT11LL_CKT W=0.34u L=40.00n
XX27 net140 DB VDD VNW PHVT11LL_CKT W=0.55u L=40.00n
XX35 net156 net171 VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX47 net172 SAN net171 VNW PHVT11LL_CKT W=0.455u L=40.00n
XX48 net172 DA VDD VNW PHVT11LL_CKT W=0.55u L=40.00n
.ENDS DXQV4_12TH40
.SUBCKT DXQV6_12TH40 CK DA DB Q SA VDD VSS
XX43 net140 SAN net171 VPW NHVT11LL_CKT W=0.21u L=40.00n
XX6 net103 c net108 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX3 net156 cn net103 VPW NHVT11LL_CKT W=0.35u L=40.00n
XX4 net104 net103 VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX9 net108 net104 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX14 net104 c net123 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX16 net124 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net123 cn net124 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 s net123 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX22 Q net123 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX26 net140 DB VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX24 SAN SA VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX34 net156 net171 VSS VPW NHVT11LL_CKT W=0.49u L=40.00n
XX45 net172 SA net171 VPW NHVT11LL_CKT W=0.21u L=40.00n
XX46 net172 DA VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX0 net156 c net103 VNW PHVT11LL_CKT W=0.25u L=40.00n
XX5 net104 net103 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX7 net103 cn net19 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net19 net104 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX15 net104 cn net123 VNW PHVT11LL_CKT W=0.445u L=40.00n
XX19 net43 s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net123 c net43 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX21 s net123 VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX23 Q net123 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX44 net140 SA net171 VNW PHVT11LL_CKT W=0.455u L=40.00n
XX25 SAN SA VDD VNW PHVT11LL_CKT W=0.34u L=40.00n
XX27 net140 DB VDD VNW PHVT11LL_CKT W=0.55u L=40.00n
XX35 net156 net171 VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX47 net172 SAN net171 VNW PHVT11LL_CKT W=0.455u L=40.00n
XX48 net172 DA VDD VNW PHVT11LL_CKT W=0.55u L=40.00n
.ENDS DXQV6_12TH40
.SUBCKT EDGRNQNV2_12TH40 CK D E QN RN VDD VSS
XX2 net0140 RN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX31 VSS net0134 net241 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net241 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net0134 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX23 m c s VPW NHVT11LL_CKT W=0.33u L=40.00n
XX21 VSS m net225 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX20 net225 c net217 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX13 net194 cn net217 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX17 m net217 VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX9 net206 s net0140 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX8 net194 en net206 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX3 net198 E net0140 VPW NHVT11LL_CKT W=0.61u L=40.00n
XX5 net194 D net198 VPW NHVT11LL_CKT W=0.46u L=40.00n
XX15 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX27 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX32 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX11 QN s VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX33 net194 RN VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX22 m cn s VNW PHVT11LL_CKT W=0.33u L=40.00n
XX12 net194 c net217 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX29 net166 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 net0134 s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX28 VDD net0134 net166 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX18 VDD m net150 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net150 cn net217 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net194 E net149 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX16 m net217 VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX6 net149 s VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net194 D net137 VNW PHVT11LL_CKT W=0.42u L=40.00n
XX0 net137 en VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX14 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX10 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX4 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX26 QN s VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
.ENDS EDGRNQNV2_12TH40
.SUBCKT EDGRNQNV4_12TH40 CK D E QN RN VDD VSS
XX2 net0140 RN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX31 VSS net0134 net241 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net241 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net0134 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX23 m c s VPW NHVT11LL_CKT W=0.33u L=40.00n
XX21 VSS m net225 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX20 net225 c net217 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX13 net194 cn net217 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX17 m net217 VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX9 net206 s net0140 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX8 net194 en net206 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX3 net198 E net0140 VPW NHVT11LL_CKT W=0.61u L=40.00n
XX5 net194 D net198 VPW NHVT11LL_CKT W=0.46u L=40.00n
XX15 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX27 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX32 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX11 QN s VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX33 net194 RN VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX22 m cn s VNW PHVT11LL_CKT W=0.42u L=40.00n
XX12 net194 c net217 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX29 net166 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 net0134 s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX28 VDD net0134 net166 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX18 VDD m net150 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net150 cn net217 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net194 E net149 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX16 m net217 VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX6 net149 s VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net194 D net137 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX0 net137 en VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX14 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX10 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX4 cn CK VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX26 QN s VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS EDGRNQNV4_12TH40
.SUBCKT EDGRNQNV6_12TH40 CK D E QN RN VDD VSS
XX2 net0140 RN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX31 VSS net0134 net241 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net241 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net0134 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX23 m c s VPW NHVT11LL_CKT W=0.33u L=40.00n
XX21 VSS m net225 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX20 net225 c net217 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX13 net194 cn net217 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX17 m net217 VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX9 net206 s net0140 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX8 net194 en net206 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX3 net198 E net0140 VPW NHVT11LL_CKT W=0.61u L=40.00n
XX5 net194 D net198 VPW NHVT11LL_CKT W=0.46u L=40.00n
XX15 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX27 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX32 cn CK VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX11 QN s VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX33 net194 RN VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX22 m cn s VNW PHVT11LL_CKT W=0.47u L=40.00n
XX12 net194 c net217 VNW PHVT11LL_CKT W=0.42u L=40.00n
XX29 net166 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 net0134 s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX28 VDD net0134 net166 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX18 VDD m net150 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net150 cn net217 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net194 E net149 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX16 m net217 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX6 net149 s VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net194 D net137 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net137 en VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX14 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX10 c cn VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX4 cn CK VDD VNW PHVT11LL_CKT W=0.16u L=40.00n
XX26 QN s VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS EDGRNQNV6_12TH40
.SUBCKT EDGRNQV2_12TH40 CK D E Q RN VDD VSS
XX2 net0140 RN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX31 VSS net0134 net241 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net241 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net0134 s VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX23 m c s VPW NHVT11LL_CKT W=0.33u L=40.00n
XX21 VSS m net225 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX20 net225 c net217 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX13 net194 cn net217 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX17 m net217 VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX9 net206 s net0140 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX8 net194 en net206 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX3 net198 E net0140 VPW NHVT11LL_CKT W=0.61u L=40.00n
XX5 net194 D net198 VPW NHVT11LL_CKT W=0.45u L=40.00n
XX15 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX27 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX32 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX11 Q net0134 VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX33 net194 RN VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX22 m cn s VNW PHVT11LL_CKT W=0.36u L=40.00n
XX12 net194 c net217 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX29 net166 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 net0134 s VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX28 VDD net0134 net166 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX18 VDD m net150 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net150 cn net217 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net194 E net149 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX16 m net217 VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX6 net149 s VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net194 D net137 VNW PHVT11LL_CKT W=0.4u L=40.00n
XX0 net137 en VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX14 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX10 c cn VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX4 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX26 Q net0134 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
.ENDS EDGRNQV2_12TH40
.SUBCKT EDGRNQV4_12TH40 CK D E Q RN VDD VSS
XX2 net0140 RN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX31 VSS net0134 net241 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net241 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net0134 s VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX23 m c s VPW NHVT11LL_CKT W=0.33u L=40.00n
XX21 VSS m net225 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX20 net225 c net217 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX13 net194 cn net217 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX17 m net217 VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX9 net206 s net0140 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX8 net194 en net206 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX3 net198 E net0140 VPW NHVT11LL_CKT W=0.61u L=40.00n
XX5 net194 D net198 VPW NHVT11LL_CKT W=0.45u L=40.00n
XX15 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX27 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX32 cn CK VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX11 Q net0134 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX33 net194 RN VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX22 m cn s VNW PHVT11LL_CKT W=0.36u L=40.00n
XX12 net194 c net217 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX29 net166 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 net0134 s VDD VNW PHVT11LL_CKT W=0.51u L=40.00n
XX28 VDD net0134 net166 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX18 VDD m net150 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net150 cn net217 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net194 E net149 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX16 m net217 VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX6 net149 s VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net194 D net137 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX0 net137 en VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX14 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX10 c cn VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX4 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX26 Q net0134 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS EDGRNQV4_12TH40
.SUBCKT EDGRNQV6_12TH40 CK D E Q RN VDD VSS
XX2 net0140 RN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX31 VSS net0134 net241 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net241 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net0134 s VSS VPW NHVT11LL_CKT W=0.37u L=40.00n
XX23 m c s VPW NHVT11LL_CKT W=0.35u L=40.00n
XX21 VSS m net225 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX20 net225 c net217 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX13 net194 cn net217 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX17 m net217 VSS VPW NHVT11LL_CKT W=0.475u L=40.00n
XX9 net206 s net0140 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX8 net194 en net206 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX3 net198 E net0140 VPW NHVT11LL_CKT W=0.61u L=40.00n
XX5 net194 D net198 VPW NHVT11LL_CKT W=0.55u L=40.00n
XX15 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX27 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX32 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX11 Q net0134 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX33 net194 RN VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX22 m cn s VNW PHVT11LL_CKT W=0.36u L=40.00n
XX12 net194 c net217 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX29 net166 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 net0134 s VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX28 VDD net0134 net166 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX18 VDD m net150 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net150 cn net217 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net194 E net149 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX16 m net217 VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX6 net149 s VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net194 D net137 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net137 en VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX14 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX10 c cn VDD VNW PHVT11LL_CKT W=0.37u L=40.00n
XX4 cn CK VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX26 Q net0134 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS EDGRNQV6_12TH40
.SUBCKT EDQNV2_12TH40 CK D E QN VDD VSS
XX31 VSS net0134 net241 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net241 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net0134 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX23 m c s VPW NHVT11LL_CKT W=0.33u L=40.00n
XX21 VSS m net225 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX20 net225 c net217 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX13 net194 cn net217 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX17 m net217 VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX9 net206 s VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX8 net194 en net206 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX3 net198 E VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX5 net194 D net198 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX15 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX27 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX32 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX11 QN s VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX22 m cn s VNW PHVT11LL_CKT W=0.33u L=40.00n
XX12 net194 c net217 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX29 net166 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 net0134 s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX28 VDD net0134 net166 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX18 VDD m net150 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net150 cn net217 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net194 E net149 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX16 m net217 VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX6 net149 s VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net194 D net137 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX0 net137 en VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX14 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX10 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX4 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX26 QN s VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
.ENDS EDQNV2_12TH40
.SUBCKT EDQNV4_12TH40 CK D E QN VDD VSS
XX31 VSS net0134 net241 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net241 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net0134 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX23 m c s VPW NHVT11LL_CKT W=0.33u L=40.00n
XX21 VSS m net225 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX20 net225 c net217 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX13 net194 cn net217 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX17 m net217 VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX9 net206 s VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX8 net194 en net206 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX3 net198 E VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX5 net194 D net198 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX15 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX27 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX32 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX11 QN s VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX22 m cn s VNW PHVT11LL_CKT W=0.36u L=40.00n
XX12 net194 c net217 VNW PHVT11LL_CKT W=0.42u L=40.00n
XX29 net166 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 net0134 s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX28 VDD net0134 net166 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX18 VDD m net150 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net150 cn net217 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net194 E net149 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX16 m net217 VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX6 net149 s VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net194 D net137 VNW PHVT11LL_CKT W=0.54u L=40.00n
XX0 net137 en VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX14 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX10 c cn VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX4 cn CK VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX26 QN s VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS EDQNV4_12TH40
.SUBCKT EDQNV6_12TH40 CK D E QN VDD VSS
XX31 VSS net0134 net241 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net241 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net0134 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX23 m c s VPW NHVT11LL_CKT W=0.33u L=40.00n
XX21 VSS m net225 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX20 net225 c net217 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX13 net194 cn net217 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX17 m net217 VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX9 net206 s VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX8 net194 en net206 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX3 net198 E VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX5 net194 D net198 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX15 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX27 c cn VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX32 cn CK VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX11 QN s VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX22 m cn s VNW PHVT11LL_CKT W=0.45u L=40.00n
XX12 net194 c net217 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX29 net166 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 net0134 s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX28 VDD net0134 net166 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX18 VDD m net150 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net150 cn net217 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net194 E net149 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX16 m net217 VDD VNW PHVT11LL_CKT W=0.59u L=40.00n
XX6 net149 s VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net194 D net137 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net137 en VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX14 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX10 c cn VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX4 cn CK VDD VNW PHVT11LL_CKT W=0.18u L=40.00n
XX26 QN s VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS EDQNV6_12TH40
.SUBCKT EDQV2_12TH40 CK D E Q VDD VSS
XX31 VSS net230 net241 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net241 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net230 s VSS VPW NHVT11LL_CKT W=0.26u L=40.00n
XX23 m c s VPW NHVT11LL_CKT W=0.26u L=40.00n
XX21 VSS m net225 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX20 net225 c net217 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX13 net194 cn net217 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX17 m net217 VSS VPW NHVT11LL_CKT W=0.46u L=40.00n
XX9 net206 s VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX8 net194 en net206 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX3 net198 E VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX5 net194 D net198 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX15 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX27 c cn VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX32 cn CK VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX11 Q net230 VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX22 m cn s VNW PHVT11LL_CKT W=0.305u L=40.00n
XX12 net194 c net217 VNW PHVT11LL_CKT W=0.28u L=40.00n
XX29 net166 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 net230 s VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX28 VDD net230 net166 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX18 VDD m net150 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net150 cn net217 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net194 E net149 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX16 m net217 VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
XX6 net149 s VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net194 D net137 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX0 net137 en VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX14 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX10 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX4 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX26 Q net230 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
.ENDS EDQV2_12TH40
.SUBCKT EDQV4_12TH40 CK D E Q VDD VSS
XX31 VSS net230 net241 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net241 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net230 s VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX23 m c s VPW NHVT11LL_CKT W=0.29u L=40.00n
XX21 VSS m net225 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX20 net225 c net217 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX13 net194 cn net217 VPW NHVT11LL_CKT W=0.26u L=40.00n
XX17 m net217 VSS VPW NHVT11LL_CKT W=0.46u L=40.00n
XX9 net206 s VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX8 net194 en net206 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX3 net198 E VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX5 net194 D net198 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX15 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX27 c cn VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX32 cn CK VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX11 Q net230 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX22 m cn s VNW PHVT11LL_CKT W=0.33u L=40.00n
XX12 net194 c net217 VNW PHVT11LL_CKT W=0.26u L=40.00n
XX29 net166 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 net230 s VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX28 VDD net230 net166 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX18 VDD m net150 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net150 cn net217 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net194 E net149 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX16 m net217 VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
XX6 net149 s VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net194 D net137 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX0 net137 en VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX14 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX10 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX4 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX26 Q net230 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS EDQV4_12TH40
.SUBCKT EDQV6_12TH40 CK D E Q VDD VSS
XX31 VSS net230 net241 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net241 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net230 s VSS VPW NHVT11LL_CKT W=0.39u L=40.00n
XX23 m c s VPW NHVT11LL_CKT W=0.36u L=40.00n
XX21 VSS m net225 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX20 net225 c net217 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX13 net194 cn net217 VPW NHVT11LL_CKT W=0.26u L=40.00n
XX17 m net217 VSS VPW NHVT11LL_CKT W=0.45u L=40.00n
XX9 net206 s VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX8 net194 en net206 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX3 net198 E VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX5 net194 D net198 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX15 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX27 c cn VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX32 cn CK VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX11 Q net230 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX22 m cn s VNW PHVT11LL_CKT W=0.41u L=40.00n
XX12 net194 c net217 VNW PHVT11LL_CKT W=0.28u L=40.00n
XX29 net166 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 net230 s VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX28 VDD net230 net166 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX18 VDD m net150 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net150 cn net217 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net194 E net149 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX16 m net217 VDD VNW PHVT11LL_CKT W=0.49u L=40.00n
XX6 net149 s VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net194 D net137 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net137 en VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX14 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX10 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX4 cn CK VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX26 Q net230 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS EDQV6_12TH40
.SUBCKT EDRNQNV2_12TH40 CK D E QN RDN VDD VSS
XX36 R RDN VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX32 net110 cn net97 VPW NHVT11LL_CKT W=330.00n L=40.00n
XX31 net110 EN net102 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net102 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX0 net106 E VSS VPW NHVT11LL_CKT W=0.59u L=40.00n
XX2 net110 D net106 VPW NHVT11LL_CKT W=0.32u L=40.00n
XX25 net122 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX27 s R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net122 net97 VSS VPW NHVT11LL_CKT W=360.00n L=40.00n
XX6 net97 c net130 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net130 net122 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net122 c s VPW NHVT11LL_CKT W=0.24u L=40.00n
XX16 net138 net140 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 s cn net138 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net140 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN s VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX35 EN E VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX37 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX33 net110 c net97 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX3 net41 EN VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX28 net37 s VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX29 net110 E net37 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net110 D net41 VNW PHVT11LL_CKT W=0.49u L=40.00n
XX26 net69 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX24 net53 R VDD VNW PHVT11LL_CKT W=0.92u L=40.00n
XX5 net122 net97 net53 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX7 net97 cn net57 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net57 net122 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net122 cn s VNW PHVT11LL_CKT W=0.37u L=40.00n
XX19 net73 net140 net69 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 s c net73 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net140 s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN s VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX34 EN E VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
.ENDS EDRNQNV2_12TH40
.SUBCKT EDRNQNV4_12TH40 CK D E QN RDN VDD VSS
XX36 R RDN VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX32 net110 cn net97 VPW NHVT11LL_CKT W=330.00n L=40.00n
XX31 net110 EN net102 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net102 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX0 net106 E VSS VPW NHVT11LL_CKT W=0.59u L=40.00n
XX2 net110 D net106 VPW NHVT11LL_CKT W=0.32u L=40.00n
XX25 net122 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX27 s R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net122 net97 VSS VPW NHVT11LL_CKT W=360.00n L=40.00n
XX6 net97 c net130 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net130 net122 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net122 c s VPW NHVT11LL_CKT W=0.24u L=40.00n
XX16 net138 net140 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 s cn net138 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net140 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN s VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX35 EN E VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX37 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX33 net110 c net97 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX3 net41 EN VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX28 net37 s VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX29 net110 E net37 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net110 D net41 VNW PHVT11LL_CKT W=0.49u L=40.00n
XX26 net69 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX24 net53 R VDD VNW PHVT11LL_CKT W=0.92u L=40.00n
XX5 net122 net97 net53 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX7 net97 cn net57 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net57 net122 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net122 cn s VNW PHVT11LL_CKT W=0.45u L=40.00n
XX19 net73 net140 net69 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 s c net73 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net140 s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN s VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX34 EN E VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.16u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.3u L=40.00n
.ENDS EDRNQNV4_12TH40
.SUBCKT EDRNQNV6_12TH40 CK D E QN RDN VDD VSS
XX36 R RDN VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX32 net110 cn net97 VPW NHVT11LL_CKT W=330.00n L=40.00n
XX31 net110 EN net102 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net102 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX0 net106 E VSS VPW NHVT11LL_CKT W=0.59u L=40.00n
XX2 net110 D net106 VPW NHVT11LL_CKT W=0.32u L=40.00n
XX25 net122 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX27 s R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net122 net97 VSS VPW NHVT11LL_CKT W=0.475u L=40.00n
XX6 net97 c net130 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net130 net122 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net122 c s VPW NHVT11LL_CKT W=0.24u L=40.00n
XX16 net138 net140 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 s cn net138 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net140 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN s VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX35 EN E VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.24u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX37 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX33 net110 c net97 VNW PHVT11LL_CKT W=0.37u L=40.00n
XX3 net41 EN VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX28 net37 s VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX29 net110 E net37 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net110 D net41 VNW PHVT11LL_CKT W=0.495u L=40.00n
XX26 net69 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX24 net53 R VDD VNW PHVT11LL_CKT W=0.92u L=40.00n
XX5 net122 net97 net53 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX7 net97 cn net57 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net57 net122 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net122 cn s VNW PHVT11LL_CKT W=0.46u L=40.00n
XX19 net73 net140 net69 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 s c net73 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net140 s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN s VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX34 EN E VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.18u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
.ENDS EDRNQNV6_12TH40
.SUBCKT EDRNQV2_12TH40 CK D E Q RDN VDD VSS
XX36 R RDN VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX32 net110 cn net97 VPW NHVT11LL_CKT W=0.26u L=40.00n
XX31 net110 EN net102 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net102 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX0 net106 E VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX2 net110 D net106 VPW NHVT11LL_CKT W=0.35u L=40.00n
XX25 net122 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX27 s R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net122 net97 VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX6 net97 c net130 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net130 net122 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net122 c s VPW NHVT11LL_CKT W=0.26u L=40.00n
XX16 net138 net140 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 s cn net138 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net140 s VSS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX22 Q net140 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX35 EN E VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX37 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX33 net110 c net97 VNW PHVT11LL_CKT W=0.31u L=40.00n
XX3 net41 EN VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX28 net37 s VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX29 net110 E net37 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net110 D net41 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX26 net69 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX24 net53 R VDD VNW PHVT11LL_CKT W=0.92u L=40.00n
XX5 net122 net97 net53 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX7 net97 cn net57 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net57 net122 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net122 cn s VNW PHVT11LL_CKT W=0.3u L=40.00n
XX19 net73 net140 net69 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 s c net73 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net140 s VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX23 Q net140 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX34 EN E VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.13u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.3u L=40.00n
.ENDS EDRNQV2_12TH40
.SUBCKT EDRNQV4_12TH40 CK D E Q RDN VDD VSS
XX36 R RDN VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX32 net110 cn net97 VPW NHVT11LL_CKT W=0.26u L=40.00n
XX31 net110 EN net102 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net102 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX0 net106 E VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX2 net110 D net106 VPW NHVT11LL_CKT W=0.35u L=40.00n
XX25 net122 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX27 s R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net122 net97 VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX6 net97 c net130 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net130 net122 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net122 c s VPW NHVT11LL_CKT W=0.26u L=40.00n
XX16 net138 net140 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 s cn net138 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net140 s VSS VPW NHVT11LL_CKT W=0.37u L=40.00n
XX22 Q net140 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX35 EN E VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX37 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX33 net110 c net97 VNW PHVT11LL_CKT W=0.31u L=40.00n
XX3 net41 EN VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX28 net37 s VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX29 net110 E net37 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net110 D net41 VNW PHVT11LL_CKT W=0.54u L=40.00n
XX26 net69 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX24 net53 R VDD VNW PHVT11LL_CKT W=0.92u L=40.00n
XX5 net122 net97 net53 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX7 net97 cn net57 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net57 net122 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net122 cn s VNW PHVT11LL_CKT W=0.3u L=40.00n
XX19 net73 net140 net69 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 s c net73 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net140 s VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX23 Q net140 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX34 EN E VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.16u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.3u L=40.00n
.ENDS EDRNQV4_12TH40
.SUBCKT EDRNQV6_12TH40 CK D E Q RDN VDD VSS
XX36 R RDN VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX32 net110 cn net97 VPW NHVT11LL_CKT W=0.26u L=40.00n
XX31 net110 EN net102 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net102 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX0 net106 E VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX2 net110 D net106 VPW NHVT11LL_CKT W=0.35u L=40.00n
XX25 net122 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX27 s R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net122 net97 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX6 net97 c net130 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net130 net122 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net122 c s VPW NHVT11LL_CKT W=0.28u L=40.00n
XX16 net138 net140 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 s cn net138 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net140 s VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX22 Q net140 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX35 EN E VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX37 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX33 net110 c net97 VNW PHVT11LL_CKT W=0.31u L=40.00n
XX3 net41 EN VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX28 net37 s VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX29 net110 E net37 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net110 D net41 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX26 net69 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX24 net53 R VDD VNW PHVT11LL_CKT W=0.92u L=40.00n
XX5 net122 net97 net53 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX7 net97 cn net57 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net57 net122 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net122 cn s VNW PHVT11LL_CKT W=0.3u L=40.00n
XX19 net73 net140 net69 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 s c net73 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net140 s VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX23 Q net140 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX34 EN E VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.16u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.3u L=40.00n
.ENDS EDRNQV6_12TH40
.SUBCKT FDCAP128_12TH40 VDD VSS
XX47 net139 net140 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX46 net143 net144 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX45 net147 net148 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX44 net151 net152 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX43 net155 net156 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX42 net159 net160 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX41 net163 net164 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX40 net167 net168 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX39 net171 net172 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX38 net175 net176 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX37 net179 net180 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX36 net183 net184 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX35 net187 net188 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX34 net191 net192 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX33 net195 net196 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX32 net199 net200 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX11 net203 net204 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX10 net207 net208 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX9 net211 net212 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX8 net215 net216 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX2 net219 net220 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX1 net223 net224 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX6 net227 net228 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX7 net231 net232 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX24 net235 net236 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX25 net239 net240 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX26 net243 net244 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX27 net247 net248 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX28 net251 net252 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX29 net255 net256 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX30 net259 net260 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX31 net263 net264 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX63 VSS net139 net140 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX62 VSS net143 net144 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX61 VSS net147 net148 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX60 VSS net151 net152 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX59 VSS net155 net156 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX58 VSS net159 net160 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX57 VSS net163 net164 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX56 VSS net167 net168 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX55 VSS net171 net172 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX54 VSS net175 net176 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX53 VSS net179 net180 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX52 VSS net183 net184 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX51 VSS net187 net188 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX50 VSS net191 net192 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX49 VSS net195 net196 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX48 VSS net199 net200 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX15 VSS net203 net204 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX14 VSS net207 net208 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX13 VSS net211 net212 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX12 VSS net215 net216 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX20 VSS net251 net252 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX19 VSS net247 net248 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX18 VSS net243 net244 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX17 VSS net239 net240 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX16 VSS net235 net236 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX5 VSS net231 net232 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX4 VSS net227 net228 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX0 VSS net223 net224 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX3 VSS net219 net220 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX23 VSS net263 net264 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX22 VSS net259 net260 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX21 VSS net255 net256 VPW NHVT11LL_CKT W=465.00n L=315.00n
.ENDS FDCAP128_12TH40
.SUBCKT FDCAP16_12TH40 VDD VSS
XX5 VSS net011 net012 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX4 VSS net015 net016 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX0 VSS net019 net020 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX3 VSS net7 net8 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX7 net011 net012 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX6 net015 net016 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX1 net019 net020 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX2 net7 net8 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
.ENDS FDCAP16_12TH40
.SUBCKT FDCAP32_12TH40 VDD VSS
XX11 net43 net44 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX10 net47 net48 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX9 net51 net52 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX8 net55 net56 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX7 net71 net72 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX6 net67 net68 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX1 net63 net64 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX2 net59 net60 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX15 VSS net43 net44 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX14 VSS net47 net48 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX13 VSS net51 net52 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX12 VSS net55 net56 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX5 VSS net71 net72 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX4 VSS net67 net68 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX0 VSS net63 net64 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX3 VSS net59 net60 VPW NHVT11LL_CKT W=465.00n L=315.00n
.ENDS FDCAP32_12TH40
.SUBCKT FDCAP4_12TH40 VDD VSS
XX3 VSS net7 net8 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX2 net7 net8 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
.ENDS FDCAP4_12TH40
.SUBCKT FDCAP64_12TH40 VDD VSS
XX23 VSS net11 net12 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX22 VSS net15 net16 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX21 VSS net19 net20 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX20 VSS net23 net24 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX19 VSS net27 net28 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX18 VSS net31 net32 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX17 VSS net35 net36 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX16 VSS net39 net40 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX12 VSS net59 net60 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX3 VSS net55 net56 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX0 VSS net51 net52 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX4 VSS net47 net48 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX5 VSS net43 net44 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX15 VSS net71 net72 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX14 VSS net67 net68 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX13 VSS net63 net64 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX31 net11 net12 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX30 net15 net16 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX29 net19 net20 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX28 net23 net24 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX27 net27 net28 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX26 net31 net32 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX25 net35 net36 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX24 net39 net40 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX11 net71 net72 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX10 net67 net68 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX9 net63 net64 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX8 net59 net60 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX2 net55 net56 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX1 net51 net52 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX6 net47 net48 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX7 net43 net44 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
.ENDS FDCAP64_12TH40
.SUBCKT FDCAP8_12TH40 VDD VSS
XX0 VSS net011 net012 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX3 VSS net7 net8 VPW NHVT11LL_CKT W=465.00n L=315.00n
XX1 net011 net012 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
XX2 net7 net8 VDD VNW PHVT11LL_CKT W=465.00n L=315.00n
.ENDS FDCAP8_12TH40
.SUBCKT FILLTIE128_12TH40 VDD VSS
.ENDS FILLTIE128_12TH40
.SUBCKT FILLTIE16_12TH40 VDD VSS
.ENDS FILLTIE16_12TH40
.SUBCKT FILLTIE32_12TH40 VDD VSS
.ENDS FILLTIE32_12TH40
.SUBCKT FILLTIE3_12TH40 VDD VSS
.ENDS FILLTIE3_12TH40
.SUBCKT FILLTIE4_12TH40 VDD VSS
.ENDS FILLTIE4_12TH40
.SUBCKT FILLTIE64_12TH40 VDD VSS
.ENDS FILLTIE64_12TH40
.SUBCKT FILLTIE8_12TH40 VDD VSS
.ENDS FILLTIE8_12TH40
.SUBCKT F_DIODE2_12TH40 A VDD VSS
DD1 A VNW PDIO11LLHVT PJ=2.9 AREA=0.1403p
DD0 VPW A NDIO11LLHVT PJ=2.9 AREA=0.1403p
.ENDS F_DIODE2_12TH40
.SUBCKT F_DIODE4_12TH40 A VDD VSS
DD1 A VNW PDIO11LLHVT PJ=5.9 AREA=0.3111p
DD0 VPW A NDIO11LLHVT PJ=5.9 AREA=0.3111p
.ENDS F_DIODE4_12TH40
.SUBCKT F_DIODE8_12TH40 A VDD VSS
DD1 A VNW PDIO11LLHVT PJ=11.9 AREA=0.6527p
DD0 VPW A NDIO11LLHVT PJ=11.9 AREA=0.6527p
.ENDS F_DIODE8_12TH40
.SUBCKT F_FILL128_12TH40 VDD VSS
.ENDS F_FILL128_12TH40
.SUBCKT F_FILL16_12TH40 VDD VSS
.ENDS F_FILL16_12TH40
.SUBCKT F_FILL1_12TH40 VDD VSS
.ENDS F_FILL1_12TH40
.SUBCKT F_FILL2_12TH40 VDD VSS
.ENDS F_FILL2_12TH40
.SUBCKT F_FILL32_12TH40 VDD VSS
.ENDS F_FILL32_12TH40
.SUBCKT F_FILL4_12TH40 VDD VSS
.ENDS F_FILL4_12TH40
.SUBCKT F_FILL64_12TH40 VDD VSS
.ENDS F_FILL64_12TH40
.SUBCKT F_FILL8_12TH40 VDD VSS
.ENDS F_FILL8_12TH40
.SUBCKT INV0SR_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=310.00n L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=270.00n L=40.00n
.ENDS INV0SR_12TH40
.SUBCKT INV0_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
.ENDS INV0_12TH40
.SUBCKT INV10SR_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=3.05u L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=2.7u L=40.00n
.ENDS INV10SR_12TH40
.SUBCKT INV10_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=2.7u L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=3.05u L=40.00n
.ENDS INV10_12TH40
.SUBCKT INV12SR_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=3.66u L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=3.24u L=40.00n
.ENDS INV12SR_12TH40
.SUBCKT INV12_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=3.24u L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
.ENDS INV12_12TH40
.SUBCKT INV16SR_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=4.88u L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=4.32u L=40.00n
.ENDS INV16SR_12TH40
.SUBCKT INV16_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=4.32u L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
.ENDS INV16_12TH40
.SUBCKT INV1SR_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=430.00n L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=380.00n L=40.00n
.ENDS INV1SR_12TH40
.SUBCKT INV1_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
.ENDS INV1_12TH40
.SUBCKT INV20SR_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=6.1u L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=5.4u L=40.00n
.ENDS INV20SR_12TH40
.SUBCKT INV20_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=5.4u L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=6.1u L=40.00n
.ENDS INV20_12TH40
.SUBCKT INV24SR_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=7.32u L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=6.48u L=40.00n
.ENDS INV24SR_12TH40
.SUBCKT INV24_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=6.48u L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=7.32u L=40.00n
.ENDS INV24_12TH40
.SUBCKT INV2SR_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
.ENDS INV2SR_12TH40
.SUBCKT INV2_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS INV2_12TH40
.SUBCKT INV32SR_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=9.76u L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=8.64u L=40.00n
.ENDS INV32SR_12TH40
.SUBCKT INV32_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=8.64u L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=9.76u L=40.00n
.ENDS INV32_12TH40
.SUBCKT INV3SR_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=860.00n L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=760.00n L=40.00n
.ENDS INV3SR_12TH40
.SUBCKT INV3_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
.ENDS INV3_12TH40
.SUBCKT INV4SR_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
.ENDS INV4SR_12TH40
.SUBCKT INV4_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS INV4_12TH40
.SUBCKT INV5SR_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=1.53u L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=1.35u L=40.00n
.ENDS INV5SR_12TH40
.SUBCKT INV5_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=1.35u L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=1.53u L=40.00n
.ENDS INV5_12TH40
.SUBCKT INV6SR_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=1.83u L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=1.62u L=40.00n
.ENDS INV6SR_12TH40
.SUBCKT INV6_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS INV6_12TH40
.SUBCKT INV7SR_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=1.88u L=40.00n
.ENDS INV7SR_12TH40
.SUBCKT INV7_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=1.88u L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
.ENDS INV7_12TH40
.SUBCKT INV8SR_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
.ENDS INV8SR_12TH40
.SUBCKT INV8_12TH40 I ZN VDD VSS
XX0 ZN I VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX3 ZN I VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS INV8_12TH40
.SUBCKT LAHQNV0_12TH40 D E QN VDD VSS
XX10 EN E VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX4 net67 net52 VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX2 net45 D VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX3 net45 E net52 VPW NHVT11LL_CKT W=0.165u L=40.00n
XX15 QN net67 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX6 net52 EN net65 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net65 net67 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX11 EN E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX5 net67 net52 VDD VNW PHVT11LL_CKT W=0.19u L=40.00n
XX1 net45 D VDD VNW PHVT11LL_CKT W=0.39u L=40.00n
XX0 net45 EN net52 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX14 QN net67 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX7 net52 E net32 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net32 net67 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS LAHQNV0_12TH40
.SUBCKT LAHQNV2_12TH40 D E QN VDD VSS
XX10 EN E VSS VPW NHVT11LL_CKT W=150.00n L=40.00n
XX4 net67 net52 VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX2 net45 D VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX3 net45 E net52 VPW NHVT11LL_CKT W=215.00n L=40.00n
XX15 QN net67 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX6 net52 EN net65 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net65 net67 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX11 EN E VDD VNW PHVT11LL_CKT W=150.00n L=40.00n
XX5 net67 net52 VDD VNW PHVT11LL_CKT W=320.00n L=40.00n
XX1 net45 D VDD VNW PHVT11LL_CKT W=480.00n L=40.00n
XX0 net45 EN net52 VNW PHVT11LL_CKT W=260.00n L=40.00n
XX14 QN net67 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX7 net52 E net32 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net32 net67 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS LAHQNV2_12TH40
.SUBCKT LAHQNV4_12TH40 D E QN VDD VSS
XX10 EN E VSS VPW NHVT11LL_CKT W=0.165u L=40.00n
XX4 net67 net52 VSS VPW NHVT11LL_CKT W=0.53u L=40.00n
XX2 net45 D VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX3 net45 E net52 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX15 QN net67 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX6 net52 EN net65 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net65 net67 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX11 EN E VDD VNW PHVT11LL_CKT W=0.165u L=40.00n
XX5 net67 net52 VDD VNW PHVT11LL_CKT W=0.53u L=40.00n
XX1 net45 D VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX0 net45 EN net52 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX14 QN net67 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX7 net52 E net32 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net32 net67 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS LAHQNV4_12TH40
.SUBCKT LAHQNV6_12TH40 D E QN VDD VSS
XX10 EN E VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX4 net67 net52 VSS VPW NHVT11LL_CKT W=0.56u L=40.00n
XX2 net45 D VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX3 net45 E net52 VPW NHVT11LL_CKT W=0.31u L=40.00n
XX15 QN net67 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX6 net52 EN net65 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net65 net67 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX11 EN E VDD VNW PHVT11LL_CKT W=0.18u L=40.00n
XX5 net67 net52 VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX1 net45 D VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX0 net45 EN net52 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX14 QN net67 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX7 net52 E net32 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net32 net67 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS LAHQNV6_12TH40
.SUBCKT LAHQNV8_12TH40 D E QN VDD VSS
XX10 EN E VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX4 net67 net52 VSS VPW NHVT11LL_CKT W=0.75u L=40.00n
XX2 net45 D VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX3 net45 E net52 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX15 QN net67 VSS VPW NHVT11LL_CKT W=2.14u L=40.00n
XX6 net52 EN net65 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net65 net67 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX11 EN E VDD VNW PHVT11LL_CKT W=0.19u L=40.00n
XX5 net67 net52 VDD VNW PHVT11LL_CKT W=0.75u L=40.00n
XX1 net45 D VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net45 EN net52 VNW PHVT11LL_CKT W=0.49u L=40.00n
XX14 QN net67 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX7 net52 E net32 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net32 net67 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS LAHQNV8_12TH40
.SUBCKT LAHQV0_12TH40 D E Q VDD VSS
XX9 net8 net28 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net19 EN net8 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX15 Q net19 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX3 net20 E net19 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX2 net20 D VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX10 EN E VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX4 net28 net19 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX8 net43 net28 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net19 E net43 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX14 Q net19 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX0 net20 EN net19 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX1 net20 D VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX11 EN E VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX5 net28 net19 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS LAHQV0_12TH40
.SUBCKT LAHQV2_12TH40 D E Q VDD VSS
XX9 net8 net28 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net19 EN net8 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX15 Q net19 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX3 net20 E net19 VPW NHVT11LL_CKT W=330.00n L=40.00n
XX2 net20 D VSS VPW NHVT11LL_CKT W=460.00n L=40.00n
XX10 EN E VSS VPW NHVT11LL_CKT W=170.00n L=40.00n
XX4 net28 net19 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX8 net43 net28 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net19 E net43 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX14 Q net19 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX0 net20 EN net19 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX1 net20 D VDD VNW PHVT11LL_CKT W=560.00n L=40.00n
XX11 EN E VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX5 net28 net19 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS LAHQV2_12TH40
.SUBCKT LAHQV4_12TH40 D E Q VDD VSS
XX9 net8 net28 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net19 EN net8 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX15 Q net19 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX3 net20 E net19 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX2 net20 D VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX10 EN E VSS VPW NHVT11LL_CKT W=170.00n L=40.00n
XX4 net28 net19 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX8 net43 net28 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net19 E net43 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX14 Q net19 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 net20 EN net19 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX1 net20 D VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX11 EN E VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX5 net28 net19 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS LAHQV4_12TH40
.SUBCKT LAHQV6_12TH40 D E Q VDD VSS
XX9 net8 net28 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net19 EN net8 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX15 Q net19 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX3 net20 E net19 VPW NHVT11LL_CKT W=0.49u L=40.00n
XX2 net20 D VSS VPW NHVT11LL_CKT W=0.56u L=40.00n
XX10 EN E VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX4 net28 net19 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX8 net43 net28 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net19 E net43 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX14 Q net19 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX0 net20 EN net19 VNW PHVT11LL_CKT W=0.49u L=40.00n
XX1 net20 D VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX11 EN E VDD VNW PHVT11LL_CKT W=0.18u L=40.00n
XX5 net28 net19 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS LAHQV6_12TH40
.SUBCKT LAHRNQNV0_12TH40 D E QN RDN VDD VSS
XX16 R RDN VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX10 EN E VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX9 net9 net13 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net13 net20 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX3 net21 E net20 VPW NHVT11LL_CKT W=0.165u L=40.00n
XX2 net21 D VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX6 net20 EN net9 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX13 net13 R VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX15 QN net13 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX17 R RDN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX11 EN E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX8 net48 net13 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net20 E net48 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net13 net20 net52 VNW PHVT11LL_CKT W=0.305u L=40.00n
XX0 net21 EN net20 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX1 net21 D VDD VNW PHVT11LL_CKT W=0.39u L=40.00n
XX14 QN net13 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX12 net52 R VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
.ENDS LAHRNQNV0_12TH40
.SUBCKT LAHRNQNV2_12TH40 D E QN RDN VDD VSS
XX16 R RDN VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX10 EN E VSS VPW NHVT11LL_CKT W=150.00n L=40.00n
XX9 net9 net13 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net13 net20 VSS VPW NHVT11LL_CKT W=180.00n L=40.00n
XX3 net21 E net20 VPW NHVT11LL_CKT W=215.00n L=40.00n
XX2 net21 D VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX6 net20 EN net9 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX13 net13 R VSS VPW NHVT11LL_CKT W=180.00n L=40.00n
XX15 QN net13 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX17 R RDN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX11 EN E VDD VNW PHVT11LL_CKT W=150.00n L=40.00n
XX8 net48 net13 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net20 E net48 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net13 net20 net52 VNW PHVT11LL_CKT W=310.00n L=40.00n
XX0 net21 EN net20 VNW PHVT11LL_CKT W=260.00n L=40.00n
XX1 net21 D VDD VNW PHVT11LL_CKT W=480.00n L=40.00n
XX14 QN net13 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX12 net52 R VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
.ENDS LAHRNQNV2_12TH40
.SUBCKT LAHRNQNV4_12TH40 D E QN RDN VDD VSS
XX16 R RDN VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX10 EN E VSS VPW NHVT11LL_CKT W=0.165u L=40.00n
XX9 net9 net13 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net13 net20 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX3 net21 E net20 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX2 net21 D VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX6 net20 EN net9 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX13 net13 R VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX15 QN net13 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX17 R RDN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX11 EN E VDD VNW PHVT11LL_CKT W=0.165u L=40.00n
XX8 net48 net13 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net20 E net48 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net13 net20 net52 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX0 net21 EN net20 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX1 net21 D VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX14 QN net13 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX12 net52 R VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
.ENDS LAHRNQNV4_12TH40
.SUBCKT LAHRNQNV6_12TH40 D E QN RDN VDD VSS
XX16 R RDN VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX10 EN E VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX9 net9 net13 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net13 net20 VSS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX3 net21 E net20 VPW NHVT11LL_CKT W=0.31u L=40.00n
XX2 net21 D VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX6 net20 EN net9 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX13 net13 R VSS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX15 QN net13 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX17 R RDN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX11 EN E VDD VNW PHVT11LL_CKT W=0.18u L=40.00n
XX8 net48 net13 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net20 E net48 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net13 net20 net52 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net21 EN net20 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX1 net21 D VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX14 QN net13 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX12 net52 R VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
.ENDS LAHRNQNV6_12TH40
.SUBCKT LAHRNQNV8_12TH40 D E QN RDN VDD VSS
XX16 R RDN VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX10 EN E VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX9 net9 net13 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net13 net20 VSS VPW NHVT11LL_CKT W=0.75u L=40.00n
XX3 net21 E net20 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX2 net21 D VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX6 net20 EN net9 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX13 net13 R VSS VPW NHVT11LL_CKT W=0.75u L=40.00n
XX15 QN net13 VSS VPW NHVT11LL_CKT W=2.14u L=40.00n
XX17 R RDN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX11 EN E VDD VNW PHVT11LL_CKT W=0.19u L=40.00n
XX8 net48 net13 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net20 E net48 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net13 net20 net52 VNW PHVT11LL_CKT W=0.62u L=40.00n
XX0 net21 EN net20 VNW PHVT11LL_CKT W=0.49u L=40.00n
XX1 net21 D VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX14 QN net13 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX12 net52 R VDD VNW PHVT11LL_CKT W=0.62u L=40.00n
.ENDS LAHRNQNV8_12TH40
.SUBCKT LAHRNQV0_12TH40 D E Q RDN VDD VSS
XX15 Q net56 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX6 net56 EN net45 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX9 net45 net57 net69 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX2 net49 D net65 VPW NHVT11LL_CKT W=0.32u L=40.00n
XX3 net49 E net56 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX4 net57 net56 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 EN E VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX16 net65 RDN VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX18 net69 RDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX14 Q net56 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX7 net56 E net12 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net12 net57 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX1 net49 D VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX0 net49 EN net56 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX5 net57 net56 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 EN E VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX17 net56 RDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS LAHRNQV0_12TH40
.SUBCKT LAHRNQV2_12TH40 D E Q RDN VDD VSS
XX15 Q net56 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX6 net56 EN net45 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX9 net45 net57 net69 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX2 net49 D net65 VPW NHVT11LL_CKT W=570.00n L=40.00n
XX3 net49 E net56 VPW NHVT11LL_CKT W=330.00n L=40.00n
XX4 net57 net56 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 EN E VSS VPW NHVT11LL_CKT W=170.00n L=40.00n
XX16 net65 RDN VSS VPW NHVT11LL_CKT W=570.00n L=40.00n
XX18 net69 RDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX14 Q net56 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX7 net56 E net12 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net12 net57 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX1 net49 D VDD VNW PHVT11LL_CKT W=445.00n L=40.00n
XX0 net49 EN net56 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX5 net57 net56 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 EN E VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX17 net56 RDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS LAHRNQV2_12TH40
.SUBCKT LAHRNQV4_12TH40 D E Q RDN VDD VSS
XX15 Q net56 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX6 net56 EN net45 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX9 net45 net57 net69 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX2 net49 D net65 VPW NHVT11LL_CKT W=570.00n L=40.00n
XX3 net49 E net56 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX4 net57 net56 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 EN E VSS VPW NHVT11LL_CKT W=170.00n L=40.00n
XX16 net65 RDN VSS VPW NHVT11LL_CKT W=570.00n L=40.00n
XX18 net69 RDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX14 Q net56 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX7 net56 E net12 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net12 net57 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX1 net49 D VDD VNW PHVT11LL_CKT W=445.00n L=40.00n
XX0 net49 EN net56 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX5 net57 net56 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 EN E VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX17 net56 RDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS LAHRNQV4_12TH40
.SUBCKT LAHRNQV6_12TH40 D E Q RDN VDD VSS
XX15 Q net56 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX6 net56 EN net45 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX9 net45 net57 net69 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX2 net49 D net65 VPW NHVT11LL_CKT W=0.61u L=40.00n
XX3 net49 E net56 VPW NHVT11LL_CKT W=0.49u L=40.00n
XX4 net57 net56 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 EN E VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX16 net65 RDN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX18 net69 RDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX14 Q net56 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX7 net56 E net12 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net12 net57 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX1 net49 D VDD VNW PHVT11LL_CKT W=0.475u L=40.00n
XX0 net49 EN net56 VNW PHVT11LL_CKT W=0.49u L=40.00n
XX5 net57 net56 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 EN E VDD VNW PHVT11LL_CKT W=0.18u L=40.00n
XX17 net56 RDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS LAHRNQV6_12TH40
.SUBCKT LAHRSNQNV2_12TH40 D E QN RDN SDN VDD VSS
XX12 net114 E net055 VPW NHVT11LL_CKT W=0.305u L=40.00n
XX6 net114 EN net99 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net107 net114 net119 VPW NHVT11LL_CKT W=0.27u L=40.00n
XX10 EN E VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX9 net99 net107 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 R RDN VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX22 QN net107 VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX27 net107 R net119 VPW NHVT11LL_CKT W=0.14u L=40.00n
XX26 net119 SDN VSS VPW NHVT11LL_CKT W=0.46u L=40.00n
XX2 net055 D VSS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX13 net114 EN net115 VNW PHVT11LL_CKT W=0.28u L=40.00n
XX25 net150 R VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX24 net107 SDN VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX1 net115 D VDD VNW PHVT11LL_CKT W=0.28u L=40.00n
XX5 net107 net114 net150 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX7 net114 E net146 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net146 net107 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 EN E VDD VNW PHVT11LL_CKT W=0.18u L=40.00n
XX23 QN net107 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX34 R RDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
.ENDS LAHRSNQNV2_12TH40
.SUBCKT LAHRSNQNV4_12TH40 D E QN RDN SDN VDD VSS
XX13 net127 EN net90 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX1 net90 D VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX11 EN E VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX25 net70 R VDD VNW PHVT11LL_CKT W=0.545u L=40.00n
XX24 net111 SDN VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX5 net111 net127 net70 VNW PHVT11LL_CKT W=0.545u L=40.00n
XX7 net127 E net66 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net66 net111 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net111 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX34 R RDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX12 net127 E net123 VPW NHVT11LL_CKT W=0.365u L=40.00n
XX2 net123 D VSS VPW NHVT11LL_CKT W=0.39u L=40.00n
XX10 EN E VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX6 net127 EN net107 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net111 net127 net91 VPW NHVT11LL_CKT W=0.32u L=40.00n
XX9 net107 net111 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 R RDN VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX22 QN net111 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX27 net111 R net91 VPW NHVT11LL_CKT W=0.14u L=40.00n
XX26 net91 SDN VSS VPW NHVT11LL_CKT W=0.46u L=40.00n
.ENDS LAHRSNQNV4_12TH40
.SUBCKT LAHRSNQNV6_12TH40 D E QN RDN SDN VDD VSS
XX13 net127 EN net90 VNW PHVT11LL_CKT W=0.4u L=40.00n
XX1 net90 D VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX11 EN E VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX25 net70 R VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX24 net111 SDN VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX5 net111 net127 net70 VNW PHVT11LL_CKT W=0.545u L=40.00n
XX7 net127 E net66 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net66 net111 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net111 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX34 R RDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX12 net127 E net123 VPW NHVT11LL_CKT W=0.435u L=40.00n
XX2 net123 D VSS VPW NHVT11LL_CKT W=0.46u L=40.00n
XX10 EN E VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX6 net127 EN net107 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net111 net127 net91 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX9 net107 net111 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 R RDN VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX22 QN net111 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX27 net111 R net91 VPW NHVT11LL_CKT W=0.14u L=40.00n
XX26 net91 SDN VSS VPW NHVT11LL_CKT W=0.46u L=40.00n
.ENDS LAHRSNQNV6_12TH40
.SUBCKT LAHRSNQV2_12TH40 D E Q RDN SDN VDD VSS
XX0 pm E net10 VPW NHVT11LL_CKT W=0.28u L=40.00n
XX1 net10 RDN net14 VPW NHVT11LL_CKT W=0.28u L=40.00n
XX2 net14 D VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX3 pm s VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX4 EN E VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX6 s SDN VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX7 Q pm VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX8 net38 pm VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX10 pm EN net46 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX11 net46 RDN net50 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX12 net50 net38 VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX13 net61 D VDD VNW PHVT11LL_CKT W=0.345u L=40.00n
XX14 net65 s net61 VNW PHVT11LL_CKT W=0.345u L=40.00n
XX15 pm EN net65 VNW PHVT11LL_CKT W=0.345u L=40.00n
XX16 net73 RDN VDD VNW PHVT11LL_CKT W=150.00n L=40.00n
XX17 pm s net73 VNW PHVT11LL_CKT W=150.00n L=40.00n
XX18 net38 pm VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX20 Q pm VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX21 s SDN VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX23 EN E VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX24 net101 net38 VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX25 net105 s net101 VNW PHVT11LL_CKT W=0.15u L=40.00n
XX26 pm E net105 VNW PHVT11LL_CKT W=0.15u L=40.00n
.ENDS LAHRSNQV2_12TH40
.SUBCKT LAHRSNQV4_12TH40 D E Q RDN SDN VDD VSS
XX0 pm E net10 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX1 net10 RDN net14 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX2 net14 D VSS VPW NHVT11LL_CKT W=0.36u L=40.00n
XX3 pm s VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX4 EN E VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX6 s SDN VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX7 Q pm VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX8 net38 pm VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX10 pm EN net46 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX11 net46 RDN net50 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX12 net50 net38 VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX13 net61 D VDD VNW PHVT11LL_CKT W=0.48u L=40.00n
XX14 net65 s net61 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX15 pm EN net65 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX16 net73 RDN VDD VNW PHVT11LL_CKT W=150.00n L=40.00n
XX17 pm s net73 VNW PHVT11LL_CKT W=150.00n L=40.00n
XX18 net38 pm VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX20 Q pm VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX21 s SDN VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX23 EN E VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX24 net101 net38 VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX25 net105 s net101 VNW PHVT11LL_CKT W=0.15u L=40.00n
XX26 pm E net105 VNW PHVT11LL_CKT W=0.15u L=40.00n
.ENDS LAHRSNQV4_12TH40
.SUBCKT LAHRSNQV6_12TH40 D E Q RDN SDN VDD VSS
XX0 net087 E net10 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX1 net10 RDN net14 VPW NHVT11LL_CKT W=0.405u L=40.00n
XX2 net14 D VSS VPW NHVT11LL_CKT W=0.405u L=40.00n
XX3 net087 s VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX4 EN E VSS VPW NHVT11LL_CKT W=0.22u L=40.00n
XX6 s SDN VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX7 Q net087 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX8 net38 net087 VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX10 net087 EN net46 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX11 net46 RDN net50 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX12 net50 net38 VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX13 net61 D VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX14 net65 s net61 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX15 net087 EN net65 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX16 net73 RDN VDD VNW PHVT11LL_CKT W=150.00n L=40.00n
XX17 net087 s net73 VNW PHVT11LL_CKT W=150.00n L=40.00n
XX18 net38 net087 VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX20 Q net087 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX21 s SDN VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX23 EN E VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX24 net101 net38 VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX25 net105 s net101 VNW PHVT11LL_CKT W=0.15u L=40.00n
XX26 net087 E net105 VNW PHVT11LL_CKT W=0.15u L=40.00n
.ENDS LAHRSNQV6_12TH40
.SUBCKT LAHSNQNV0_12TH40 D E QN SDN VDD VSS
XX10 EN E VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX4 net63 net52 net65 VPW NHVT11LL_CKT W=0.21u L=40.00n
XX2 net45 D VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX3 net45 E net52 VPW NHVT11LL_CKT W=0.165u L=40.00n
XX15 QN net63 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX6 net52 EN net61 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net61 net63 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net65 SDN VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX11 EN E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX5 net63 net52 VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX1 net45 D VDD VNW PHVT11LL_CKT W=0.39u L=40.00n
XX0 net45 EN net52 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX14 QN net63 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX7 net52 E net28 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net28 net63 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX12 net63 SDN VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
.ENDS LAHSNQNV0_12TH40
.SUBCKT LAHSNQNV2_12TH40 D E QN SDN VDD VSS
XX10 EN E VSS VPW NHVT11LL_CKT W=150.00n L=40.00n
XX4 net63 net52 net65 VPW NHVT11LL_CKT W=290.00n L=40.00n
XX2 net45 D VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX3 net45 E net52 VPW NHVT11LL_CKT W=215.00n L=40.00n
XX15 QN net63 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX6 net52 EN net61 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net61 net63 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net65 SDN VSS VPW NHVT11LL_CKT W=290.00n L=40.00n
XX11 EN E VDD VNW PHVT11LL_CKT W=150.00n L=40.00n
XX5 net63 net52 VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX1 net45 D VDD VNW PHVT11LL_CKT W=480.00n L=40.00n
XX0 net45 EN net52 VNW PHVT11LL_CKT W=260.00n L=40.00n
XX14 QN net63 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX7 net52 E net28 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net28 net63 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX12 net63 SDN VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
.ENDS LAHSNQNV2_12TH40
.SUBCKT LAHSNQNV4_12TH40 D E QN SDN VDD VSS
XX10 EN E VSS VPW NHVT11LL_CKT W=0.165u L=40.00n
XX4 net63 net52 net65 VPW NHVT11LL_CKT W=0.58u L=40.00n
XX2 net45 D VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX3 net45 E net52 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX15 QN net63 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX6 net52 EN net61 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net61 net63 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net65 SDN VSS VPW NHVT11LL_CKT W=0.58u L=40.00n
XX11 EN E VDD VNW PHVT11LL_CKT W=0.165u L=40.00n
XX5 net63 net52 VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX1 net45 D VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX0 net45 EN net52 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX14 QN net63 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX7 net52 E net28 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net28 net63 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX12 net63 SDN VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
.ENDS LAHSNQNV4_12TH40
.SUBCKT LAHSNQNV6_12TH40 D E QN SDN VDD VSS
XX10 EN E VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX4 net63 net52 net65 VPW NHVT11LL_CKT W=0.61u L=40.00n
XX2 net45 D VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX3 net45 E net52 VPW NHVT11LL_CKT W=0.31u L=40.00n
XX15 QN net63 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX6 net52 EN net61 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net61 net63 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net65 SDN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX11 EN E VDD VNW PHVT11LL_CKT W=0.18u L=40.00n
XX5 net63 net52 VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX1 net45 D VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX0 net45 EN net52 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX14 QN net63 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX7 net52 E net28 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net28 net63 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX12 net63 SDN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
.ENDS LAHSNQNV6_12TH40
.SUBCKT LAHSNQNV8_12TH40 D E QN SDN VDD VSS
XX10 EN E VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX4 net63 net52 net65 VPW NHVT11LL_CKT W=1.18u L=40.00n
XX2 net45 D VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX3 net45 E net52 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX15 QN net63 VSS VPW NHVT11LL_CKT W=2.14u L=40.00n
XX6 net52 EN net61 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net61 net63 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net65 SDN VSS VPW NHVT11LL_CKT W=1.18u L=40.00n
XX11 EN E VDD VNW PHVT11LL_CKT W=0.19u L=40.00n
XX5 net63 net52 VDD VNW PHVT11LL_CKT W=0.67u L=40.00n
XX1 net45 D VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net45 EN net52 VNW PHVT11LL_CKT W=0.49u L=40.00n
XX14 QN net63 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX7 net52 E net28 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net28 net63 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX12 net63 SDN VDD VNW PHVT11LL_CKT W=0.67u L=40.00n
.ENDS LAHSNQNV8_12TH40
.SUBCKT LAHSNQV2_12TH40 D E Q SDN VDD VSS
XX17 S SDN VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX9 net5 net7 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net28 EN net5 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX15 Q net28 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX4 net7 net28 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 EN E VSS VPW NHVT11LL_CKT W=170.00n L=40.00n
XX3 net29 E net28 VPW NHVT11LL_CKT W=220.00n L=40.00n
XX2 net29 D VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX16 net28 S VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 S SDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX12 net68 S VDD VNW PHVT11LL_CKT W=510.00n L=40.00n
XX8 net48 net7 net44 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX7 net28 E net48 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX14 Q net28 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX5 net7 net28 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 EN E VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX0 net29 EN net28 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX1 net29 D net68 VNW PHVT11LL_CKT W=510.00n L=40.00n
XX13 net44 S VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
.ENDS LAHSNQV2_12TH40
.SUBCKT LAHSNQV4_12TH40 D E Q SDN VDD VSS
XX17 S SDN VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX9 net5 net7 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net28 EN net5 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX15 Q net28 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX4 net7 net28 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 EN E VSS VPW NHVT11LL_CKT W=170.00n L=40.00n
XX3 net29 E net28 VPW NHVT11LL_CKT W=0.24u L=40.00n
XX2 net29 D VSS VPW NHVT11LL_CKT W=0.24u L=40.00n
XX16 net28 S VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 S SDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX12 net68 S VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX8 net48 net7 net44 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX7 net28 E net48 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX14 Q net28 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX5 net7 net28 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 EN E VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX0 net29 EN net28 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX1 net29 D net68 VNW PHVT11LL_CKT W=0.56u L=40.00n
XX13 net44 S VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
.ENDS LAHSNQV4_12TH40
.SUBCKT LAHSNQV6_12TH40 D E Q SDN VDD VSS
XX17 S SDN VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX9 net5 net7 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net28 EN net5 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX15 Q net28 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX4 net7 net28 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 EN E VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX3 net29 E net28 VPW NHVT11LL_CKT W=0.32u L=40.00n
XX2 net29 D VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX16 net28 S VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 S SDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX12 net68 S VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX8 net48 net7 net44 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX7 net28 E net48 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX14 Q net28 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX5 net7 net28 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 EN E VDD VNW PHVT11LL_CKT W=0.18u L=40.00n
XX0 net29 EN net28 VNW PHVT11LL_CKT W=0.49u L=40.00n
XX1 net29 D net68 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX13 net44 S VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
.ENDS LAHSNQV6_12TH40
.SUBCKT LALQNV0_12TH40 D EN QN VDD VSS
XX6 net63 EN net68 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net56 D VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX3 net56 ENN net63 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX4 net92 net63 VSS VPW NHVT11LL_CKT W=0.175u L=40.00n
XX9 net68 net92 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 ENN EN VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net92 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX1 net56 D VDD VNW PHVT11LL_CKT W=0.39u L=40.00n
XX0 net56 EN net63 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX5 net92 net63 VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX7 net63 ENN net19 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net19 net92 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 ENN EN VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
XX23 QN net92 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
.ENDS LALQNV0_12TH40
.SUBCKT LALQNV2_12TH40 D EN QN VDD VSS
XX6 net63 EN net68 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net56 D VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX3 net56 ENN net63 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX4 net92 net63 VSS VPW NHVT11LL_CKT W=300.00n L=40.00n
XX9 net68 net92 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 ENN EN VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net92 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX1 net56 D VDD VNW PHVT11LL_CKT W=480.00n L=40.00n
XX0 net56 EN net63 VNW PHVT11LL_CKT W=260.00n L=40.00n
XX5 net92 net63 VDD VNW PHVT11LL_CKT W=345.00n L=40.00n
XX7 net63 ENN net19 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net19 net92 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 ENN EN VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
XX23 QN net92 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS LALQNV2_12TH40
.SUBCKT LALQNV4_12TH40 D EN QN VDD VSS
XX6 net63 EN net68 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net56 D VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX3 net56 ENN net63 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX4 net92 net63 VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX9 net68 net92 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 ENN EN VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net92 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX1 net56 D VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX0 net56 EN net63 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX5 net92 net63 VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX7 net63 ENN net19 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net19 net92 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 ENN EN VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
XX23 QN net92 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS LALQNV4_12TH40
.SUBCKT LALQNV6_12TH40 D EN QN VDD VSS
XX6 net63 EN net68 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net56 D VSS VPW NHVT11LL_CKT W=0.49u L=40.00n
XX3 net56 ENN net63 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX4 net92 net63 VSS VPW NHVT11LL_CKT W=0.51u L=40.00n
XX9 net68 net92 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 ENN EN VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net92 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX1 net56 D VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX0 net56 EN net63 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX5 net92 net63 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX7 net63 ENN net19 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net19 net92 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 ENN EN VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
XX23 QN net92 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS LALQNV6_12TH40
.SUBCKT LALQNV8_12TH40 D EN QN VDD VSS
XX6 net63 EN net68 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net56 D VSS VPW NHVT11LL_CKT W=0.49u L=40.00n
XX3 net56 ENN net63 VPW NHVT11LL_CKT W=0.49u L=40.00n
XX4 net92 net63 VSS VPW NHVT11LL_CKT W=0.68u L=40.00n
XX9 net68 net92 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 ENN EN VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net92 VSS VPW NHVT11LL_CKT W=2.14u L=40.00n
XX1 net56 D VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX0 net56 EN net63 VNW PHVT11LL_CKT W=0.49u L=40.00n
XX5 net92 net63 VDD VNW PHVT11LL_CKT W=0.82u L=40.00n
XX7 net63 ENN net19 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net19 net92 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 ENN EN VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
XX23 QN net92 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS LALQNV8_12TH40
.SUBCKT LALQV0_12TH40 D EN Q VDD VSS
XX10 ENN EN VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net12 net16 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net16 net23 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX3 net24 ENN net23 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX2 net24 D VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX6 net23 EN net12 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 Q net23 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX11 ENN EN VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
XX8 net47 net16 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net23 ENN net47 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net16 net23 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX0 net24 EN net23 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX1 net24 D VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX23 Q net23 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
.ENDS LALQV0_12TH40
.SUBCKT LALQV2_12TH40 D EN Q VDD VSS
XX10 ENN EN VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net12 net16 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net16 net23 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX3 net24 ENN net23 VPW NHVT11LL_CKT W=330.00n L=40.00n
XX2 net24 D VSS VPW NHVT11LL_CKT W=475.00n L=40.00n
XX6 net23 EN net12 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 Q net23 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX11 ENN EN VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
XX8 net47 net16 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net23 ENN net47 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net16 net23 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX0 net24 EN net23 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX1 net24 D VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX23 Q net23 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS LALQV2_12TH40
.SUBCKT LALQV4_12TH40 D EN Q VDD VSS
XX10 ENN EN VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net12 net16 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net16 net23 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX3 net24 ENN net23 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX2 net24 D VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX6 net23 EN net12 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 Q net23 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX11 ENN EN VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
XX8 net47 net16 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net23 ENN net47 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net16 net23 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX0 net24 EN net23 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX1 net24 D VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX23 Q net23 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS LALQV4_12TH40
.SUBCKT LALQV6_12TH40 D EN Q VDD VSS
XX10 ENN EN VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net12 net16 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net16 net23 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX3 net24 ENN net23 VPW NHVT11LL_CKT W=0.49u L=40.00n
XX2 net24 D VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX6 net23 EN net12 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 Q net23 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX11 ENN EN VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
XX8 net47 net16 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net23 ENN net47 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net16 net23 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX0 net24 EN net23 VNW PHVT11LL_CKT W=0.49u L=40.00n
XX1 net24 D VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX23 Q net23 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS LALQV6_12TH40
.SUBCKT LALRNQNV2_12TH40 D EN QN RDN VDD VSS
XX16 R RDN VSS VPW NHVT11LL_CKT W=0.22u L=40.00n
XX15 QN net44 VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX13 net44 R VSS VPW NHVT11LL_CKT W=180.00n L=40.00n
XX6 net43 EN net48 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net36 D VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX3 net36 ENN net43 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX4 net44 net43 VSS VPW NHVT11LL_CKT W=180.00n L=40.00n
XX9 net48 net44 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 ENN EN VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 R RDN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX12 net0129 R VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
XX14 QN net44 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 net36 D VDD VNW PHVT11LL_CKT W=480.00n L=40.00n
XX0 net36 EN net43 VNW PHVT11LL_CKT W=260.00n L=40.00n
XX5 net44 net43 net0129 VNW PHVT11LL_CKT W=310.00n L=40.00n
XX7 net43 ENN net19 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net19 net44 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 ENN EN VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
.ENDS LALRNQNV2_12TH40
.SUBCKT LALRNQNV4_12TH40 D EN QN RDN VDD VSS
XX16 R RDN VSS VPW NHVT11LL_CKT W=0.22u L=40.00n
XX15 QN net44 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX13 net44 R VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX6 net43 EN net48 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net36 D VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX3 net36 ENN net43 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX4 net44 net43 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX9 net48 net44 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 ENN EN VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 R RDN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX12 net0129 R VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX14 QN net44 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 net36 D VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX0 net36 EN net43 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX5 net44 net43 net0129 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX7 net43 ENN net19 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net19 net44 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 ENN EN VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
.ENDS LALRNQNV4_12TH40
.SUBCKT LALRNQNV6_12TH40 D EN QN RDN VDD VSS
XX16 R RDN VSS VPW NHVT11LL_CKT W=0.22u L=40.00n
XX15 QN net44 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX13 net44 R VSS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX6 net43 EN net48 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net36 D VSS VPW NHVT11LL_CKT W=0.49u L=40.00n
XX3 net36 ENN net43 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX4 net44 net43 VSS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX9 net48 net44 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 ENN EN VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 R RDN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX12 net0129 R VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX14 QN net44 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX1 net36 D VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX0 net36 EN net43 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX5 net44 net43 net0129 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX7 net43 ENN net19 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net19 net44 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 ENN EN VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
.ENDS LALRNQNV6_12TH40
.SUBCKT LALRNQV2_12TH40 D EN Q RDN VDD VSS
XX18 net13 RDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX16 net25 RDN VSS VPW NHVT11LL_CKT W=570.00n L=40.00n
XX10 ENN EN VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net9 net36 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX3 net37 ENN net36 VPW NHVT11LL_CKT W=330.00n L=40.00n
XX2 net37 D net25 VPW NHVT11LL_CKT W=570.00n L=40.00n
XX9 net17 net9 net13 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX6 net36 EN net17 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX15 Q net36 VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX17 net36 RDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 ENN EN VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
XX5 net9 net36 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX0 net37 EN net36 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX1 net37 D VDD VNW PHVT11LL_CKT W=445.00n L=40.00n
XX8 net60 net9 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net36 ENN net60 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX14 Q net36 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS LALRNQV2_12TH40
.SUBCKT LALRNQV4_12TH40 D EN Q RDN VDD VSS
XX18 net13 RDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX16 net25 RDN VSS VPW NHVT11LL_CKT W=570.00n L=40.00n
XX10 ENN EN VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net9 net36 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX3 net37 ENN net36 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX2 net37 D net25 VPW NHVT11LL_CKT W=570.00n L=40.00n
XX9 net17 net9 net13 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX6 net36 EN net17 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX15 Q net36 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX17 net36 RDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 ENN EN VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
XX5 net9 net36 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX0 net37 EN net36 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX1 net37 D VDD VNW PHVT11LL_CKT W=445.00n L=40.00n
XX8 net60 net9 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net36 ENN net60 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX14 Q net36 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS LALRNQV4_12TH40
.SUBCKT LALRNQV6_12TH40 D EN Q RDN VDD VSS
XX18 net13 RDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX16 net25 RDN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX10 ENN EN VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net9 net36 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX3 net37 ENN net36 VPW NHVT11LL_CKT W=0.49u L=40.00n
XX2 net37 D net25 VPW NHVT11LL_CKT W=0.61u L=40.00n
XX9 net17 net9 net13 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX6 net36 EN net17 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX15 Q net36 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX17 net36 RDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 ENN EN VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
XX5 net9 net36 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX0 net37 EN net36 VNW PHVT11LL_CKT W=0.49u L=40.00n
XX1 net37 D VDD VNW PHVT11LL_CKT W=0.475u L=40.00n
XX8 net60 net9 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net36 ENN net60 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX14 Q net36 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS LALRNQV6_12TH40
.SUBCKT LALRSNQNV2_12TH40 D EN QN RDN SDN VDD VSS
XX13 net69 EN net058 VNW PHVT11LL_CKT W=0.28u L=40.00n
XX1 net058 D VDD VNW PHVT11LL_CKT W=0.28u L=40.00n
XX25 net29 R VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX24 net70 SDN VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX5 net70 net69 net29 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX7 net69 ENN net33 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net33 net70 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 ENN EN VDD VNW PHVT11LL_CKT W=0.26u L=40.00n
XX23 QN net70 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX34 R RDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX2 net091 D VSS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX12 net69 ENN net091 VPW NHVT11LL_CKT W=0.305u L=40.00n
XX27 net70 R net58 VPW NHVT11LL_CKT W=0.14u L=40.00n
XX26 net58 SDN VSS VPW NHVT11LL_CKT W=0.46u L=40.00n
XX4 net70 net69 net58 VPW NHVT11LL_CKT W=0.27u L=40.00n
XX6 net69 EN net78 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net78 net70 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 ENN EN VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX22 QN net70 VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX33 R RDN VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
.ENDS LALRSNQNV2_12TH40
.SUBCKT LALRSNQNV4_12TH40 D EN QN RDN SDN VDD VSS
XX9 net59 net67 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net67 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX33 R RDN VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX2 net87 D VSS VPW NHVT11LL_CKT W=0.39u L=40.00n
XX12 net83 ENN net87 VPW NHVT11LL_CKT W=0.365u L=40.00n
XX10 ENN EN VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX27 net67 R net71 VPW NHVT11LL_CKT W=0.14u L=40.00n
XX26 net71 SDN VSS VPW NHVT11LL_CKT W=0.46u L=40.00n
XX4 net67 net83 net71 VPW NHVT11LL_CKT W=0.32u L=40.00n
XX6 net83 EN net59 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX1 net126 D VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX13 net83 EN net126 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX11 ENN EN VDD VNW PHVT11LL_CKT W=0.26u L=40.00n
XX25 net110 R VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX24 net67 SDN VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX5 net67 net83 net110 VNW PHVT11LL_CKT W=0.54u L=40.00n
XX7 net83 ENN net106 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net106 net67 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net67 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX34 R RDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
.ENDS LALRSNQNV4_12TH40
.SUBCKT LALRSNQNV6_12TH40 D EN QN RDN SDN VDD VSS
XX9 net59 net67 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net67 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX33 R RDN VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX2 net87 D VSS VPW NHVT11LL_CKT W=0.46u L=40.00n
XX12 net83 ENN net87 VPW NHVT11LL_CKT W=0.435u L=40.00n
XX10 ENN EN VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX27 net67 R net71 VPW NHVT11LL_CKT W=0.14u L=40.00n
XX26 net71 SDN VSS VPW NHVT11LL_CKT W=0.46u L=40.00n
XX4 net67 net83 net71 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX6 net83 EN net59 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX1 net126 D VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX13 net83 EN net126 VNW PHVT11LL_CKT W=0.4u L=40.00n
XX11 ENN EN VDD VNW PHVT11LL_CKT W=0.26u L=40.00n
XX25 net110 R VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX24 net67 SDN VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX5 net67 net83 net110 VNW PHVT11LL_CKT W=0.54u L=40.00n
XX7 net83 ENN net106 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net106 net67 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net67 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX34 R RDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
.ENDS LALRSNQNV6_12TH40
.SUBCKT LALRSNQV2_12TH40 D EN Q RDN SDN VDD VSS
XX1 Q pm VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX2 s SDN VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX4 ENN EN VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX5 net22 D VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX6 net26 RDN net22 VPW NHVT11LL_CKT W=0.28u L=40.00n
XX7 pm ENN net26 VPW NHVT11LL_CKT W=0.28u L=40.00n
XX8 pm s VSS VPW NHVT11LL_CKT W=140.00n L=40.00n
XX9 net38 pm VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX10 net42 net38 VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX11 net46 RDN net42 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX12 pm EN net46 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX13 net61 D VDD VNW PHVT11LL_CKT W=0.345u L=40.00n
XX14 net65 s net61 VNW PHVT11LL_CKT W=0.345u L=40.00n
XX15 pm EN net65 VNW PHVT11LL_CKT W=0.345u L=40.00n
XX16 net73 RDN VDD VNW PHVT11LL_CKT W=150.00n L=40.00n
XX17 pm s net73 VNW PHVT11LL_CKT W=150.00n L=40.00n
XX18 net38 pm VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX20 ENN EN VDD VNW PHVT11LL_CKT W=0.26u L=40.00n
XX22 s SDN VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX23 Q pm VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX24 net101 net38 VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX25 net105 s net101 VNW PHVT11LL_CKT W=0.15u L=40.00n
XX26 pm ENN net105 VNW PHVT11LL_CKT W=0.15u L=40.00n
.ENDS LALRSNQV2_12TH40
.SUBCKT LALRSNQV4_12TH40 D EN Q RDN SDN VDD VSS
XX1 Q pm VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX2 s SDN VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX4 ENN EN VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX5 net22 D VSS VPW NHVT11LL_CKT W=0.36u L=40.00n
XX6 net26 RDN net22 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX7 pm ENN net26 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX8 pm s VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX9 net38 pm VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX10 net42 net38 VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX11 net46 RDN net42 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX12 pm EN net46 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX13 net61 D VDD VNW PHVT11LL_CKT W=0.48u L=40.00n
XX14 net65 s net61 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX15 pm EN net65 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX16 net73 RDN VDD VNW PHVT11LL_CKT W=150.00n L=40.00n
XX17 pm s net73 VNW PHVT11LL_CKT W=150.00n L=40.00n
XX18 net38 pm VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX20 ENN EN VDD VNW PHVT11LL_CKT W=0.26u L=40.00n
XX22 s SDN VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX23 Q pm VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX24 net101 net38 VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX25 net105 s net101 VNW PHVT11LL_CKT W=0.15u L=40.00n
XX26 pm ENN net105 VNW PHVT11LL_CKT W=0.15u L=40.00n
.ENDS LALRSNQV4_12TH40
.SUBCKT LALRSNQV6_12TH40 D EN Q RDN SDN VDD VSS
XX1 Q pm VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX2 s SDN VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX4 ENN EN VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX5 net22 D VSS VPW NHVT11LL_CKT W=0.36u L=40.00n
XX6 net26 RDN net22 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX7 pm ENN net26 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX8 pm s VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX9 net38 pm VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX10 net42 net38 VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX11 net46 RDN net42 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX12 pm EN net46 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX13 net61 D VDD VNW PHVT11LL_CKT W=0.48u L=40.00n
XX14 net65 s net61 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX15 pm EN net65 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX16 net73 RDN VDD VNW PHVT11LL_CKT W=150.00n L=40.00n
XX17 pm s net73 VNW PHVT11LL_CKT W=150.00n L=40.00n
XX18 net38 pm VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX20 ENN EN VDD VNW PHVT11LL_CKT W=0.26u L=40.00n
XX22 s SDN VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX23 Q pm VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX24 net101 net38 VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX25 net105 s net101 VNW PHVT11LL_CKT W=0.15u L=40.00n
XX26 pm ENN net105 VNW PHVT11LL_CKT W=0.15u L=40.00n
.ENDS LALRSNQV6_12TH40
.SUBCKT LALSNQNV0_12TH40 D EN QN SDN VDD VSS
XX16 net5 SDN VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX9 net13 net15 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net24 EN net13 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX15 QN net15 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX3 net25 ENN net24 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX2 net25 D VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX4 net15 net24 net5 VPW NHVT11LL_CKT W=0.21u L=40.00n
XX10 ENN EN VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX12 net15 SDN VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX8 net52 net15 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net24 ENN net52 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX14 QN net15 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX0 net25 EN net24 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX1 net25 D VDD VNW PHVT11LL_CKT W=0.39u L=40.00n
XX5 net15 net24 VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX11 ENN EN VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
.ENDS LALSNQNV0_12TH40
.SUBCKT LALSNQNV2_12TH40 D EN QN SDN VDD VSS
XX16 net5 SDN VSS VPW NHVT11LL_CKT W=290.00n L=40.00n
XX9 net13 net15 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net24 EN net13 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX15 QN net15 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX3 net25 ENN net24 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX2 net25 D VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX4 net15 net24 net5 VPW NHVT11LL_CKT W=290.00n L=40.00n
XX10 ENN EN VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX12 net15 SDN VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX8 net52 net15 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net24 ENN net52 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX14 QN net15 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX0 net25 EN net24 VNW PHVT11LL_CKT W=260.00n L=40.00n
XX1 net25 D VDD VNW PHVT11LL_CKT W=480.00n L=40.00n
XX5 net15 net24 VDD VNW PHVT11LL_CKT W=170.00n L=40.00n
XX11 ENN EN VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
.ENDS LALSNQNV2_12TH40
.SUBCKT LALSNQNV4_12TH40 D EN QN SDN VDD VSS
XX16 net5 SDN VSS VPW NHVT11LL_CKT W=0.58u L=40.00n
XX9 net13 net15 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net24 EN net13 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX15 QN net15 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX3 net25 ENN net24 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX2 net25 D VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX4 net15 net24 net5 VPW NHVT11LL_CKT W=0.58u L=40.00n
XX10 ENN EN VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX12 net15 SDN VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX8 net52 net15 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net24 ENN net52 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX14 QN net15 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 net25 EN net24 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX1 net25 D VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX5 net15 net24 VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX11 ENN EN VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
.ENDS LALSNQNV4_12TH40
.SUBCKT LALSNQNV6_12TH40 D EN QN SDN VDD VSS
XX16 net5 SDN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX9 net13 net15 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net24 EN net13 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX15 QN net15 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX3 net25 ENN net24 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX2 net25 D VSS VPW NHVT11LL_CKT W=0.49u L=40.00n
XX4 net15 net24 net5 VPW NHVT11LL_CKT W=0.61u L=40.00n
XX10 ENN EN VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX12 net15 SDN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX8 net52 net15 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net24 ENN net52 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX14 QN net15 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX0 net25 EN net24 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX1 net25 D VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX5 net15 net24 VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX11 ENN EN VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
.ENDS LALSNQNV6_12TH40
.SUBCKT LALSNQNV8_12TH40 D EN QN SDN VDD VSS
XX16 net5 SDN VSS VPW NHVT11LL_CKT W=1.18u L=40.00n
XX9 net13 net15 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net24 EN net13 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX15 QN net15 VSS VPW NHVT11LL_CKT W=2.14u L=40.00n
XX3 net25 ENN net24 VPW NHVT11LL_CKT W=0.49u L=40.00n
XX2 net25 D VSS VPW NHVT11LL_CKT W=0.49u L=40.00n
XX4 net15 net24 net5 VPW NHVT11LL_CKT W=1.18u L=40.00n
XX10 ENN EN VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX12 net15 SDN VDD VNW PHVT11LL_CKT W=0.67u L=40.00n
XX8 net52 net15 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net24 ENN net52 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX14 QN net15 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX0 net25 EN net24 VNW PHVT11LL_CKT W=0.49u L=40.00n
XX1 net25 D VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX5 net15 net24 VDD VNW PHVT11LL_CKT W=0.67u L=40.00n
XX11 ENN EN VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
.ENDS LALSNQNV8_12TH40
.SUBCKT LALSNQV2_12TH40 D EN Q SDN VDD VSS
XX17 S SDN VSS VPW NHVT11LL_CKT W=0.22u L=40.00n
XX16 net44 S VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net37 D VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX3 net37 ENN net44 VPW NHVT11LL_CKT W=330.00n L=40.00n
XX10 ENN EN VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net53 net44 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX15 Q net44 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX6 net44 EN net65 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net65 net53 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 S SDN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX13 net0153 S VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX1 net37 D net0137 VNW PHVT11LL_CKT W=510.00n L=40.00n
XX0 net37 EN net44 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX11 ENN EN VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
XX5 net53 net44 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX14 Q net44 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX7 net44 ENN net32 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX8 net32 net53 net0153 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX12 net0137 S VDD VNW PHVT11LL_CKT W=510.00n L=40.00n
.ENDS LALSNQV2_12TH40
.SUBCKT LALSNQV4_12TH40 D EN Q SDN VDD VSS
XX17 S SDN VSS VPW NHVT11LL_CKT W=0.22u L=40.00n
XX16 net44 S VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net37 D VSS VPW NHVT11LL_CKT W=0.24u L=40.00n
XX3 net37 ENN net44 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX10 ENN EN VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net53 net44 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX15 Q net44 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX6 net44 EN net65 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net65 net53 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 S SDN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX13 net0153 S VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX1 net37 D net0137 VNW PHVT11LL_CKT W=0.56u L=40.00n
XX0 net37 EN net44 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX11 ENN EN VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
XX5 net53 net44 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX14 Q net44 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX7 net44 ENN net32 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX8 net32 net53 net0153 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX12 net0137 S VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
.ENDS LALSNQV4_12TH40
.SUBCKT LALSNQV6_12TH40 D EN Q SDN VDD VSS
XX17 S SDN VSS VPW NHVT11LL_CKT W=0.22u L=40.00n
XX16 net44 S VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net37 D VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX3 net37 ENN net44 VPW NHVT11LL_CKT W=0.46u L=40.00n
XX10 ENN EN VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net53 net44 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX15 Q net44 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX6 net44 EN net65 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net65 net53 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 S SDN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX13 net0153 S VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX1 net37 D net0137 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net37 EN net44 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX11 ENN EN VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
XX5 net53 net44 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX14 Q net44 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX7 net44 ENN net32 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX8 net32 net53 net0153 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX12 net0137 S VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
.ENDS LALSNQV6_12TH40
.SUBCKT MAJ23V2_12TH40 A1 A2 A3 Z VDD VSS
XX11 Z net33 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX4 net33 A3 net37 VPW NHVT11LL_CKT W=300.00n L=40.00n
XX2 net37 A1 VSS VPW NHVT11LL_CKT W=300.00n L=40.00n
XX5 net37 A2 VSS VPW NHVT11LL_CKT W=300.00n L=40.00n
XX8 net33 A1 net49 VPW NHVT11LL_CKT W=300.00n L=40.00n
XX9 net49 A2 VSS VPW NHVT11LL_CKT W=300.00n L=40.00n
XX1 net9 A1 VDD VNW PHVT11LL_CKT W=360.00n L=40.00n
XX0 net9 A2 VDD VNW PHVT11LL_CKT W=360.00n L=40.00n
XX3 net33 A3 net9 VNW PHVT11LL_CKT W=360.00n L=40.00n
XX6 net28 A2 VDD VNW PHVT11LL_CKT W=360.00n L=40.00n
XX7 net33 A1 net28 VNW PHVT11LL_CKT W=360.00n L=40.00n
XX10 Z net33 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS MAJ23V2_12TH40
.SUBCKT MAJ23V3_12TH40 A1 A2 A3 Z VDD VSS
XX11 Z net33 VSS VPW NHVT11LL_CKT W=0.75u L=40.00n
XX4 net33 A3 net37 VPW NHVT11LL_CKT W=0.375u L=40.00n
XX2 net37 A1 VSS VPW NHVT11LL_CKT W=0.375u L=40.00n
XX5 net37 A2 VSS VPW NHVT11LL_CKT W=0.375u L=40.00n
XX8 net33 A1 net49 VPW NHVT11LL_CKT W=0.375u L=40.00n
XX9 net49 A2 VSS VPW NHVT11LL_CKT W=0.375u L=40.00n
XX1 net9 A1 VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
XX0 net9 A2 VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
XX3 net33 A3 net9 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX6 net28 A2 VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
XX7 net33 A1 net28 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX10 Z net33 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
.ENDS MAJ23V3_12TH40
.SUBCKT MAJ23V4_12TH40 A1 A2 A3 Z VDD VSS
XX11 Z net33 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX4 net33 A3 net37 VPW NHVT11LL_CKT W=0.505u L=40.00n
XX2 net37 A1 VSS VPW NHVT11LL_CKT W=0.505u L=40.00n
XX5 net37 A2 VSS VPW NHVT11LL_CKT W=0.505u L=40.00n
XX8 net33 A1 net49 VPW NHVT11LL_CKT W=0.505u L=40.00n
XX9 net49 A2 VSS VPW NHVT11LL_CKT W=0.505u L=40.00n
XX1 net9 A1 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net9 A2 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX3 net33 A3 net9 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX6 net28 A2 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX7 net33 A1 net28 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX10 Z net33 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS MAJ23V4_12TH40
.SUBCKT MAOI222V1_12TH40 A B C ZN VDD VSS
XX9 net5 C VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX5 net9 B VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX4 net13 A VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX13 ZN B net5 VPW NHVT11LL_CKT W=270.00n L=40.00n
XX8 ZN A net9 VPW NHVT11LL_CKT W=270.00n L=40.00n
XX11 ZN C net13 VPW NHVT11LL_CKT W=270.00n L=40.00n
XX12 net44 A VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX7 net44 C VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX6 ZN A net48 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX3 net48 B net44 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX2 ZN B net48 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX10 net48 C net44 VNW PHVT11LL_CKT W=430.00n L=40.00n
.ENDS MAOI222V1_12TH40
.SUBCKT MAOI222V2_12TH40 A B C ZN VDD VSS
XX9 net5 C VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX5 net9 B VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX4 net13 A VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX13 ZN B net5 VPW NHVT11LL_CKT W=380.00n L=40.00n
XX8 ZN A net9 VPW NHVT11LL_CKT W=380.00n L=40.00n
XX11 ZN C net13 VPW NHVT11LL_CKT W=380.00n L=40.00n
XX12 net44 A VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX7 net44 C VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX6 ZN A net48 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX3 net48 B net44 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX2 ZN B net48 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX10 net48 C net44 VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS MAOI222V2_12TH40
.SUBCKT MAOI222V4_12TH40 A B C ZN VDD VSS
XX9 net5 C VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX5 net9 B VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX4 net13 A VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX13 ZN B net5 VPW NHVT11LL_CKT W=760.00n L=40.00n
XX8 ZN A net9 VPW NHVT11LL_CKT W=760.00n L=40.00n
XX11 ZN C net13 VPW NHVT11LL_CKT W=760.00n L=40.00n
XX12 net44 A VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX7 net44 C VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX6 ZN A net48 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX3 net48 B net44 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX2 ZN B net48 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX10 net48 C net44 VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS MAOI222V4_12TH40
.SUBCKT MAOI222V8_12TH40 A B C ZN VDD VSS
XX9 net5 C VSS VPW NHVT11LL_CKT W=1.52u L=40.00n
XX5 net9 B VSS VPW NHVT11LL_CKT W=1.52u L=40.00n
XX4 net13 A VSS VPW NHVT11LL_CKT W=1.52u L=40.00n
XX13 ZN B net5 VPW NHVT11LL_CKT W=1.52u L=40.00n
XX8 ZN A net9 VPW NHVT11LL_CKT W=1.52u L=40.00n
XX11 ZN C net13 VPW NHVT11LL_CKT W=1.52u L=40.00n
XX12 net44 A VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX7 net44 C VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX6 ZN A net48 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX3 net48 B net44 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX2 ZN B net48 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX10 net48 C net44 VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS MAOI222V8_12TH40
.SUBCKT MUX2NV0_12TH40 I0 I1 S ZN VDD VSS
XX10 SN S VSS VPW NHVT11LL_CKT W=0.435u L=40.00n
XX7 BN S ZN VPW NHVT11LL_CKT W=0.25u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX5 AN SN ZN VPW NHVT11LL_CKT W=0.25u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX11 SN S VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX6 BN SN ZN VNW PHVT11LL_CKT W=0.25u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX4 AN S ZN VNW PHVT11LL_CKT W=0.25u L=40.00n
.ENDS MUX2NV0_12TH40
.SUBCKT MUX2NV1_12TH40 I0 I1 S ZN VDD VSS
XX10 SN S VSS VPW NHVT11LL_CKT W=0.48u L=40.00n
XX7 BN S ZN VPW NHVT11LL_CKT W=0.35u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX5 AN SN ZN VPW NHVT11LL_CKT W=0.35u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX11 SN S VDD VNW PHVT11LL_CKT W=0.55u L=40.00n
XX6 BN SN ZN VNW PHVT11LL_CKT W=0.35u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX4 AN S ZN VNW PHVT11LL_CKT W=0.35u L=40.00n
.ENDS MUX2NV1_12TH40
.SUBCKT MUX2NV2_12TH40 I0 I1 S ZN VDD VSS
XX10 SN S VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX7 BN S ZN VPW NHVT11LL_CKT W=500.00n L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX5 AN SN ZN VPW NHVT11LL_CKT W=500.00n L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX11 SN S VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX6 BN SN ZN VNW PHVT11LL_CKT W=500.00n L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX4 AN S ZN VNW PHVT11LL_CKT W=500.00n L=40.00n
.ENDS MUX2NV2_12TH40
.SUBCKT MUX2NV3_12TH40 I0 I1 S ZN VDD VSS
XX10 SN S VSS VPW NHVT11LL_CKT W=0.79u L=40.00n
XX7 BN S ZN VPW NHVT11LL_CKT W=0.7u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=0.7u L=40.00n
XX5 AN SN ZN VPW NHVT11LL_CKT W=0.7u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=0.7u L=40.00n
XX11 SN S VDD VNW PHVT11LL_CKT W=0.9u L=40.00n
XX6 BN SN ZN VNW PHVT11LL_CKT W=0.7u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=0.8u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=0.8u L=40.00n
XX4 AN S ZN VNW PHVT11LL_CKT W=0.7u L=40.00n
.ENDS MUX2NV3_12TH40
.SUBCKT MUX2NV4_12TH40 I0 I1 S ZN VDD VSS
XX10 SN S VSS VPW NHVT11LL_CKT W=0.93u L=40.00n
XX7 BN S ZN VPW NHVT11LL_CKT W=1u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=1u L=40.00n
XX5 AN SN ZN VPW NHVT11LL_CKT W=1u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=1u L=40.00n
XX11 SN S VDD VNW PHVT11LL_CKT W=1.06u L=40.00n
XX6 BN SN ZN VNW PHVT11LL_CKT W=1u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=1.14u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=1.14u L=40.00n
XX4 AN S ZN VNW PHVT11LL_CKT W=1u L=40.00n
.ENDS MUX2NV4_12TH40
.SUBCKT MUX2NV6_12TH40 I0 I1 S ZN VDD VSS
XX10 SN S VSS VPW NHVT11LL_CKT W=1.32u L=40.00n
XX7 BN S ZN VPW NHVT11LL_CKT W=1.5u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=1.5u L=40.00n
XX5 AN SN ZN VPW NHVT11LL_CKT W=1.5u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=1.5u L=40.00n
XX11 SN S VDD VNW PHVT11LL_CKT W=1.53u L=40.00n
XX6 BN SN ZN VNW PHVT11LL_CKT W=1.5u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=1.71u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=1.71u L=40.00n
XX4 AN S ZN VNW PHVT11LL_CKT W=1.5u L=40.00n
.ENDS MUX2NV6_12TH40
.SUBCKT MUX2NV8_12TH40 I0 I1 S ZN VDD VSS
XX10 SN S VSS VPW NHVT11LL_CKT W=1.72u L=40.00n
XX7 BN S ZN VPW NHVT11LL_CKT W=2u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=2u L=40.00n
XX5 AN SN ZN VPW NHVT11LL_CKT W=2u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=2u L=40.00n
XX11 SN S VDD VNW PHVT11LL_CKT W=1.96u L=40.00n
XX6 BN SN ZN VNW PHVT11LL_CKT W=2u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=2.28u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=2.28u L=40.00n
XX4 AN S ZN VNW PHVT11LL_CKT W=2u L=40.00n
.ENDS MUX2NV8_12TH40
.SUBCKT MUX2V0_12TH40 I0 I1 S Z VDD VSS
XX7 BN S net40 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX5 AN SN net40 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX8 Z net40 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX10 SN S VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX6 BN SN net40 VNW PHVT11LL_CKT W=0.24u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=0.24u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=0.24u L=40.00n
XX4 AN S net40 VNW PHVT11LL_CKT W=0.24u L=40.00n
XX9 Z net40 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX11 SN S VDD VNW PHVT11LL_CKT W=0.24u L=40.00n
.ENDS MUX2V0_12TH40
.SUBCKT MUX2V12_12TH40 I0 I1 S Z VDD VSS
XX7 BN S net40 VPW NHVT11LL_CKT W=1.245u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=1.245u L=40.00n
XX5 AN SN net40 VPW NHVT11LL_CKT W=1.245u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=1.245u L=40.00n
XX8 Z net40 VSS VPW NHVT11LL_CKT W=3.21u L=40.00n
XX10 SN S VSS VPW NHVT11LL_CKT W=0.82u L=40.00n
XX6 BN SN net40 VNW PHVT11LL_CKT W=1.5u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=1.5u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=1.5u L=40.00n
XX4 AN S net40 VNW PHVT11LL_CKT W=1.5u L=40.00n
XX9 Z net40 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX11 SN S VDD VNW PHVT11LL_CKT W=0.93u L=40.00n
.ENDS MUX2V12_12TH40
.SUBCKT MUX2V1_12TH40 I0 I1 S Z VDD VSS
XX7 BN S net40 VPW NHVT11LL_CKT W=0.24u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=0.24u L=40.00n
XX5 AN SN net40 VPW NHVT11LL_CKT W=0.24u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=0.24u L=40.00n
XX8 Z net40 VSS VPW NHVT11LL_CKT W=0.375u L=40.00n
XX10 SN S VSS VPW NHVT11LL_CKT W=0.24u L=40.00n
XX6 BN SN net40 VNW PHVT11LL_CKT W=0.295u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=0.295u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=0.295u L=40.00n
XX4 AN S net40 VNW PHVT11LL_CKT W=0.295u L=40.00n
XX9 Z net40 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX11 SN S VDD VNW PHVT11LL_CKT W=0.27u L=40.00n
.ENDS MUX2V1_12TH40
.SUBCKT MUX2V2_12TH40 I0 I1 S Z VDD VSS
XX7 BN S net40 VPW NHVT11LL_CKT W=300.00n L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=300.00n L=40.00n
XX5 AN SN net40 VPW NHVT11LL_CKT W=300.00n L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=300.00n L=40.00n
XX8 Z net40 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX10 SN S VSS VPW NHVT11LL_CKT W=285.00n L=40.00n
XX6 BN SN net40 VNW PHVT11LL_CKT W=360.00n L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=360.00n L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=360.00n L=40.00n
XX4 AN S net40 VNW PHVT11LL_CKT W=360.00n L=40.00n
XX9 Z net40 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX11 SN S VDD VNW PHVT11LL_CKT W=325.00n L=40.00n
.ENDS MUX2V2_12TH40
.SUBCKT MUX2V3_12TH40 I0 I1 S Z VDD VSS
XX7 BN S net40 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=0.41u L=40.00n
XX5 AN SN net40 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=0.41u L=40.00n
XX8 Z net40 VSS VPW NHVT11LL_CKT W=0.75u L=40.00n
XX10 SN S VSS VPW NHVT11LL_CKT W=0.37u L=40.00n
XX6 BN SN net40 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX4 AN S net40 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX9 Z net40 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX11 SN S VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
.ENDS MUX2V3_12TH40
.SUBCKT MUX2V4_12TH40 I0 I1 S Z VDD VSS
XX7 BN S net40 VPW NHVT11LL_CKT W=0.5u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX5 AN SN net40 VPW NHVT11LL_CKT W=0.5u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX8 Z net40 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX10 SN S VSS VPW NHVT11LL_CKT W=0.41u L=40.00n
XX6 BN SN net40 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX4 AN S net40 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX9 Z net40 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX11 SN S VDD VNW PHVT11LL_CKT W=0.47u L=40.00n
.ENDS MUX2V4_12TH40
.SUBCKT MUX2V6_12TH40 I0 I1 S Z VDD VSS
XX7 BN S net40 VPW NHVT11LL_CKT W=0.76u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=0.76u L=40.00n
XX5 AN SN net40 VPW NHVT11LL_CKT W=0.76u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=0.76u L=40.00n
XX8 Z net40 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX10 SN S VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX6 BN SN net40 VNW PHVT11LL_CKT W=0.93u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=0.93u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=0.93u L=40.00n
XX4 AN S net40 VNW PHVT11LL_CKT W=0.93u L=40.00n
XX9 Z net40 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX11 SN S VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
.ENDS MUX2V6_12TH40
.SUBCKT MUX2V8_12TH40 I0 I1 S Z VDD VSS
XX7 BN S net40 VPW NHVT11LL_CKT W=0.83u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=0.83u L=40.00n
XX5 AN SN net40 VPW NHVT11LL_CKT W=0.83u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=0.83u L=40.00n
XX8 Z net40 VSS VPW NHVT11LL_CKT W=2.14u L=40.00n
XX10 SN S VSS VPW NHVT11LL_CKT W=0.58u L=40.00n
XX6 BN SN net40 VNW PHVT11LL_CKT W=1u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=1u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=1u L=40.00n
XX4 AN S net40 VNW PHVT11LL_CKT W=1u L=40.00n
XX9 Z net40 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX11 SN S VDD VNW PHVT11LL_CKT W=0.66u L=40.00n
.ENDS MUX2V8_12TH40
.SUBCKT MUX3NV1_12TH40 I0 I1 I2 S0 S1 ZN VDD VSS
XX0 net71 S1 net58 VPW NHVT11LL_CKT W=290.00n L=40.00n
XX12 net67 S1N net58 VPW NHVT11LL_CKT W=290.00n L=40.00n
XX14 ZN net58 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX22 net67 net90 VSS VPW NHVT11LL_CKT W=290.00n L=40.00n
XX21 net71 net91 VSS VPW NHVT11LL_CKT W=290.00n L=40.00n
XX3 net75 I0 VSS VPW NHVT11LL_CKT W=290.00n L=40.00n
XX4 net79 I1 VSS VPW NHVT11LL_CKT W=290.00n L=40.00n
XX9 net75 S0N net90 VPW NHVT11LL_CKT W=290.00n L=40.00n
XX10 net79 S0 net90 VPW NHVT11LL_CKT W=290.00n L=40.00n
XX1 net91 I2 VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX17 S0N S0 VSS VPW NHVT11LL_CKT W=310.00n L=40.00n
XX18 S1N S1 VSS VPW NHVT11LL_CKT W=310.00n L=40.00n
XX6 net71 S1N net58 VNW PHVT11LL_CKT W=350.00n L=40.00n
XX15 ZN net58 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX13 net67 S1 net58 VNW PHVT11LL_CKT W=350.00n L=40.00n
XX23 net67 net90 VDD VNW PHVT11LL_CKT W=350.00n L=40.00n
XX20 net71 net91 VDD VNW PHVT11LL_CKT W=350.00n L=40.00n
XX2 net75 I0 VDD VNW PHVT11LL_CKT W=350.00n L=40.00n
XX5 net79 I1 VDD VNW PHVT11LL_CKT W=350.00n L=40.00n
XX8 net75 S0 net90 VNW PHVT11LL_CKT W=350.00n L=40.00n
XX11 net79 S0N net90 VNW PHVT11LL_CKT W=350.00n L=40.00n
XX7 net91 I2 VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX16 S0N S0 VDD VNW PHVT11LL_CKT W=350.00n L=40.00n
XX19 S1N S1 VDD VNW PHVT11LL_CKT W=350.00n L=40.00n
.ENDS MUX3NV1_12TH40
.SUBCKT MUX3NV2_12TH40 I0 I1 I2 S0 S1 ZN VDD VSS
XX0 net71 S1 net58 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX12 net67 S1N net58 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX14 ZN net58 VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX22 net67 net90 VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX21 net71 net91 VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX3 net75 I0 VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX4 net79 I1 VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX9 net75 S0N net90 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX10 net79 S0 net90 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX1 net91 I2 VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX17 S0N S0 VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX18 S1N S1 VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX6 net71 S1N net58 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX15 ZN net58 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX13 net67 S1 net58 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX23 net67 net90 VDD VNW PHVT11LL_CKT W=390.00n L=40.00n
XX20 net71 net91 VDD VNW PHVT11LL_CKT W=390.00n L=40.00n
XX2 net75 I0 VDD VNW PHVT11LL_CKT W=390.00n L=40.00n
XX5 net79 I1 VDD VNW PHVT11LL_CKT W=390.00n L=40.00n
XX8 net75 S0 net90 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX11 net79 S0N net90 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX7 net91 I2 VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX16 S0N S0 VDD VNW PHVT11LL_CKT W=370.00n L=40.00n
XX19 S1N S1 VDD VNW PHVT11LL_CKT W=370.00n L=40.00n
.ENDS MUX3NV2_12TH40
.SUBCKT MUX3NV4_12TH40 I0 I1 I2 S0 S1 ZN VDD VSS
XX0 net71 S1 net58 VPW NHVT11LL_CKT W=380.00n L=40.00n
XX12 net67 S1N net58 VPW NHVT11LL_CKT W=380.00n L=40.00n
XX14 ZN net58 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX22 net67 net90 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX21 net71 net91 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX3 net75 I0 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX4 net79 I1 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX9 net75 S0N net90 VPW NHVT11LL_CKT W=380.00n L=40.00n
XX10 net79 S0 net90 VPW NHVT11LL_CKT W=380.00n L=40.00n
XX1 net91 I2 VSS VPW NHVT11LL_CKT W=240.00n L=40.00n
XX17 S0N S0 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX18 S1N S1 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX6 net71 S1N net58 VNW PHVT11LL_CKT W=460.00n L=40.00n
XX15 ZN net58 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX13 net67 S1 net58 VNW PHVT11LL_CKT W=460.00n L=40.00n
XX23 net67 net90 VDD VNW PHVT11LL_CKT W=460.00n L=40.00n
XX20 net71 net91 VDD VNW PHVT11LL_CKT W=460.00n L=40.00n
XX2 net75 I0 VDD VNW PHVT11LL_CKT W=460.00n L=40.00n
XX5 net79 I1 VDD VNW PHVT11LL_CKT W=460.00n L=40.00n
XX8 net75 S0 net90 VNW PHVT11LL_CKT W=460.00n L=40.00n
XX11 net79 S0N net90 VNW PHVT11LL_CKT W=460.00n L=40.00n
XX7 net91 I2 VDD VNW PHVT11LL_CKT W=300.00n L=40.00n
XX16 S0N S0 VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX19 S1N S1 VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
.ENDS MUX3NV4_12TH40
.SUBCKT MUX3NV8_12TH40 I0 I1 I2 S0 S1 ZN VDD VSS
XX0 net71 S1 net58 VPW NHVT11LL_CKT W=970.00n L=40.00n
XX12 net67 S1N net58 VPW NHVT11LL_CKT W=970.00n L=40.00n
XX14 ZN net58 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX22 net67 net90 VSS VPW NHVT11LL_CKT W=970.00n L=40.00n
XX21 net71 net91 VSS VPW NHVT11LL_CKT W=970.00n L=40.00n
XX3 net75 I0 VSS VPW NHVT11LL_CKT W=970.00n L=40.00n
XX4 net79 I1 VSS VPW NHVT11LL_CKT W=970.00n L=40.00n
XX9 net75 S0N net90 VPW NHVT11LL_CKT W=970.00n L=40.00n
XX10 net79 S0 net90 VPW NHVT11LL_CKT W=970.00n L=40.00n
XX1 net91 I2 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX17 S0N S0 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX18 S1N S1 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX6 net71 S1N net58 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX15 ZN net58 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX13 net67 S1 net58 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX23 net67 net90 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX20 net71 net91 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX2 net75 I0 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX5 net79 I1 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX8 net75 S0 net90 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX11 net79 S0N net90 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX7 net91 I2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX16 S0N S0 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX19 S1N S1 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS MUX3NV8_12TH40
.SUBCKT MUX3V1_12TH40 I0 I1 I2 S0 S1 Z VDD VSS
XX18 S1N S1 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX17 S0N S0 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX14 Z net30 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX12 net34 S1N net30 VPW NHVT11LL_CKT W=280.00n L=40.00n
XX1 net23 I2 VSS VPW NHVT11LL_CKT W=280.00n L=40.00n
XX0 net23 S1 net30 VPW NHVT11LL_CKT W=280.00n L=40.00n
XX10 net39 S0 net34 VPW NHVT11LL_CKT W=280.00n L=40.00n
XX9 net43 S0N net34 VPW NHVT11LL_CKT W=280.00n L=40.00n
XX4 net39 I1 VSS VPW NHVT11LL_CKT W=280.00n L=40.00n
XX3 net43 I0 VSS VPW NHVT11LL_CKT W=280.00n L=40.00n
XX19 S1N S1 VDD VNW PHVT11LL_CKT W=290.00n L=40.00n
XX16 S0N S0 VDD VNW PHVT11LL_CKT W=290.00n L=40.00n
XX13 net34 S1 net30 VNW PHVT11LL_CKT W=350.00n L=40.00n
XX15 Z net30 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX7 net23 I2 VDD VNW PHVT11LL_CKT W=350.00n L=40.00n
XX6 net23 S1N net30 VNW PHVT11LL_CKT W=350.00n L=40.00n
XX11 net39 S0N net34 VNW PHVT11LL_CKT W=0.35u L=40.00n
XX8 net43 S0 net34 VNW PHVT11LL_CKT W=350.00n L=40.00n
XX5 net39 I1 VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX2 net43 I0 VDD VNW PHVT11LL_CKT W=350.00n L=40.00n
.ENDS MUX3V1_12TH40
.SUBCKT MUX3V2_12TH40 I0 I1 I2 S0 S1 Z VDD VSS
XX18 S1N S1 VSS VPW NHVT11LL_CKT W=280.00n L=40.00n
XX17 S0N S0 VSS VPW NHVT11LL_CKT W=280.00n L=40.00n
XX14 Z net30 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX12 net34 S1N net30 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX1 net23 I2 VSS VPW NHVT11LL_CKT W=340.00n L=40.00n
XX0 net23 S1 net30 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX10 net39 S0 net34 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX9 net43 S0N net34 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX4 net39 I1 VSS VPW NHVT11LL_CKT W=340.00n L=40.00n
XX3 net43 I0 VSS VPW NHVT11LL_CKT W=340.00n L=40.00n
XX19 S1N S1 VDD VNW PHVT11LL_CKT W=320.00n L=40.00n
XX16 S0N S0 VDD VNW PHVT11LL_CKT W=320.00n L=40.00n
XX13 net34 S1 net30 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX15 Z net30 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX7 net23 I2 VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX6 net23 S1N net30 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX11 net39 S0N net34 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX8 net43 S0 net34 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX5 net39 I1 VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX2 net43 I0 VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
.ENDS MUX3V2_12TH40
.SUBCKT MUX3V4_12TH40 I0 I1 I2 S0 S1 Z VDD VSS
XX18 S1N S1 VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX17 S0N S0 VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX14 Z net30 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX12 net34 S1N net30 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX1 net23 I2 VSS VPW NHVT11LL_CKT W=690.00n L=40.00n
XX0 net23 S1 net30 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX10 net39 S0 net34 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX9 net43 S0N net34 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX4 net39 I1 VSS VPW NHVT11LL_CKT W=690.00n L=40.00n
XX3 net43 I0 VSS VPW NHVT11LL_CKT W=690.00n L=40.00n
XX19 S1N S1 VDD VNW PHVT11LL_CKT W=580.00n L=40.00n
XX16 S0N S0 VDD VNW PHVT11LL_CKT W=580.00n L=40.00n
XX13 net34 S1 net30 VNW PHVT11LL_CKT W=870.00n L=40.00n
XX15 Z net30 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX7 net23 I2 VDD VNW PHVT11LL_CKT W=870.00n L=40.00n
XX6 net23 S1N net30 VNW PHVT11LL_CKT W=870.00n L=40.00n
XX11 net39 S0N net34 VNW PHVT11LL_CKT W=870.00n L=40.00n
XX8 net43 S0 net34 VNW PHVT11LL_CKT W=870.00n L=40.00n
XX5 net39 I1 VDD VNW PHVT11LL_CKT W=870.00n L=40.00n
XX2 net43 I0 VDD VNW PHVT11LL_CKT W=870.00n L=40.00n
.ENDS MUX3V4_12TH40
.SUBCKT MUX3V8_12TH40 I0 I1 I2 S0 S1 Z VDD VSS
XX18 S1N S1 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX17 S0N S0 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX14 Z net30 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX12 net34 S1N net30 VPW NHVT11LL_CKT W=970.00n L=40.00n
XX1 net23 I2 VSS VPW NHVT11LL_CKT W=970.00n L=40.00n
XX0 net23 S1 net30 VPW NHVT11LL_CKT W=970.00n L=40.00n
XX10 net39 S0 net34 VPW NHVT11LL_CKT W=970.00n L=40.00n
XX9 net43 S0N net34 VPW NHVT11LL_CKT W=970.00n L=40.00n
XX4 net39 I1 VSS VPW NHVT11LL_CKT W=970.00n L=40.00n
XX3 net43 I0 VSS VPW NHVT11LL_CKT W=970.00n L=40.00n
XX19 S1N S1 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX16 S0N S0 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX13 net34 S1 net30 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX15 Z net30 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX7 net23 I2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX6 net23 S1N net30 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX11 net39 S0N net34 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX8 net43 S0 net34 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX5 net39 I1 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX2 net43 I0 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS MUX3V8_12TH40
.SUBCKT MUX4NV0_12TH40 I0 I1 I2 I3 S0 S1 ZN VDD VSS
XX29 S0N S0 VSS VPW NHVT11LL_CKT W=0.42u L=40.00n
XX26 S1N S1 VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX24 ZN net23 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX22 net48 S1N net23 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX20 net44 S1 net23 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX14 DN S0 net35 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX13 CN S0N net35 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX12 CN I2 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX11 DN I3 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX10 net44 net35 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX5 AN S0N net63 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX7 BN S0 net63 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX8 net48 net63 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX28 S0N S0 VDD VNW PHVT11LL_CKT W=0.48u L=40.00n
XX27 S1N S1 VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX25 ZN net23 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX23 net48 S1 net23 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX21 net44 S1N net23 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX19 DN S0N net35 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX18 CN S0 net35 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX17 CN I2 VDD VNW PHVT11LL_CKT W=0.3u L=40.00n
XX16 DN I3 VDD VNW PHVT11LL_CKT W=0.3u L=40.00n
XX15 net44 net35 VDD VNW PHVT11LL_CKT W=0.3u L=40.00n
XX9 net48 net63 VDD VNW PHVT11LL_CKT W=0.3u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=0.3u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=0.3u L=40.00n
XX4 AN S0 net63 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX6 BN S0N net63 VNW PHVT11LL_CKT W=0.3u L=40.00n
.ENDS MUX4NV0_12TH40
.SUBCKT MUX4NV1_12TH40 I0 I1 I2 I3 S0 S1 ZN VDD VSS
XX29 S0N S0 VSS VPW NHVT11LL_CKT W=0.46u L=40.00n
XX26 S1N S1 VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX24 ZN net23 VSS VPW NHVT11LL_CKT W=0.375u L=40.00n
XX22 net48 S1N net23 VPW NHVT11LL_CKT W=0.29u L=40.00n
XX20 net44 S1 net23 VPW NHVT11LL_CKT W=0.29u L=40.00n
XX14 DN S0 net35 VPW NHVT11LL_CKT W=0.29u L=40.00n
XX13 CN S0N net35 VPW NHVT11LL_CKT W=0.29u L=40.00n
XX12 CN I2 VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX11 DN I3 VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX10 net44 net35 VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX5 AN S0N net63 VPW NHVT11LL_CKT W=0.29u L=40.00n
XX7 BN S0 net63 VPW NHVT11LL_CKT W=0.29u L=40.00n
XX8 net48 net63 VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX28 S0N S0 VDD VNW PHVT11LL_CKT W=0.53u L=40.00n
XX27 S1N S1 VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX25 ZN net23 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX23 net48 S1 net23 VNW PHVT11LL_CKT W=0.35u L=40.00n
XX21 net44 S1N net23 VNW PHVT11LL_CKT W=0.35u L=40.00n
XX19 DN S0N net35 VNW PHVT11LL_CKT W=0.35u L=40.00n
XX18 CN S0 net35 VNW PHVT11LL_CKT W=0.35u L=40.00n
XX17 CN I2 VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX16 DN I3 VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX15 net44 net35 VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX9 net48 net63 VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX4 AN S0 net63 VNW PHVT11LL_CKT W=0.35u L=40.00n
XX6 BN S0N net63 VNW PHVT11LL_CKT W=0.35u L=40.00n
.ENDS MUX4NV1_12TH40
.SUBCKT MUX4NV2_12TH40 I0 I1 I2 I3 S0 S1 ZN VDD VSS
XX29 S0N S0 VSS VPW NHVT11LL_CKT W=495.00n L=40.00n
XX26 S1N S1 VSS VPW NHVT11LL_CKT W=325.00n L=40.00n
XX24 ZN net23 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX22 net48 S1N net23 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX20 net44 S1 net23 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX14 DN S0 net35 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX13 CN S0N net35 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX12 CN I2 VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX11 DN I3 VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX10 net44 net35 VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX5 AN S0N net63 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX7 BN S0 net63 VPW NHVT11LL_CKT W=320.00n L=40.00n
XX8 net48 net63 VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX28 S0N S0 VDD VNW PHVT11LL_CKT W=565.00n L=40.00n
XX27 S1N S1 VDD VNW PHVT11LL_CKT W=370.00n L=40.00n
XX25 ZN net23 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX23 net48 S1 net23 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX21 net44 S1N net23 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX19 DN S0N net35 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX18 CN S0 net35 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX17 CN I2 VDD VNW PHVT11LL_CKT W=390.00n L=40.00n
XX16 DN I3 VDD VNW PHVT11LL_CKT W=390.00n L=40.00n
XX15 net44 net35 VDD VNW PHVT11LL_CKT W=390.00n L=40.00n
XX9 net48 net63 VDD VNW PHVT11LL_CKT W=390.00n L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=390.00n L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=390.00n L=40.00n
XX4 AN S0 net63 VNW PHVT11LL_CKT W=390.00n L=40.00n
XX6 BN S0N net63 VNW PHVT11LL_CKT W=390.00n L=40.00n
.ENDS MUX4NV2_12TH40
.SUBCKT MUX4NV3_12TH40 I0 I1 I2 I3 S0 S1 ZN VDD VSS
XX29 S0N S0 VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX26 S1N S1 VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX24 ZN net23 VSS VPW NHVT11LL_CKT W=0.75u L=40.00n
XX22 net48 S1N net23 VPW NHVT11LL_CKT W=0.35u L=40.00n
XX20 net44 S1 net23 VPW NHVT11LL_CKT W=0.35u L=40.00n
XX14 DN S0 net35 VPW NHVT11LL_CKT W=0.35u L=40.00n
XX13 CN S0N net35 VPW NHVT11LL_CKT W=0.35u L=40.00n
XX12 CN I2 VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX11 DN I3 VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX10 net44 net35 VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX5 AN S0N net63 VPW NHVT11LL_CKT W=0.35u L=40.00n
XX7 BN S0 net63 VPW NHVT11LL_CKT W=0.35u L=40.00n
XX8 net48 net63 VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX28 S0N S0 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX27 S1N S1 VDD VNW PHVT11LL_CKT W=0.39u L=40.00n
XX25 ZN net23 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX23 net48 S1 net23 VNW PHVT11LL_CKT W=0.425u L=40.00n
XX21 net44 S1N net23 VNW PHVT11LL_CKT W=0.425u L=40.00n
XX19 DN S0N net35 VNW PHVT11LL_CKT W=0.425u L=40.00n
XX18 CN S0 net35 VNW PHVT11LL_CKT W=0.425u L=40.00n
XX17 CN I2 VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX16 DN I3 VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX15 net44 net35 VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX9 net48 net63 VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX4 AN S0 net63 VNW PHVT11LL_CKT W=0.425u L=40.00n
XX6 BN S0N net63 VNW PHVT11LL_CKT W=0.425u L=40.00n
.ENDS MUX4NV3_12TH40
.SUBCKT MUX4NV4_12TH40 I0 I1 I2 I3 S0 S1 ZN VDD VSS
XX29 S0N S0 VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX26 S1N S1 VSS VPW NHVT11LL_CKT W=0.355u L=40.00n
XX24 ZN net23 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX22 net48 S1N net23 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX20 net44 S1 net23 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX14 DN S0 net35 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX13 CN S0N net35 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX12 CN I2 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX11 DN I3 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX10 net44 net35 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX5 AN S0N net63 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX7 BN S0 net63 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX8 net48 net63 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX28 S0N S0 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX27 S1N S1 VDD VNW PHVT11LL_CKT W=0.405u L=40.00n
XX25 ZN net23 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX23 net48 S1 net23 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX21 net44 S1N net23 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX19 DN S0N net35 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX18 CN S0 net35 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX17 CN I2 VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
XX16 DN I3 VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
XX15 net44 net35 VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
XX9 net48 net63 VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
XX4 AN S0 net63 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX6 BN S0N net63 VNW PHVT11LL_CKT W=0.46u L=40.00n
.ENDS MUX4NV4_12TH40
.SUBCKT MUX4NV6_12TH40 I0 I1 I2 I3 S0 S1 ZN VDD VSS
XX29 S0N S0 VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX26 S1N S1 VSS VPW NHVT11LL_CKT W=0.37u L=40.00n
XX24 ZN net23 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX22 net48 S1N net23 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX20 net44 S1 net23 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX14 DN S0 net35 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX13 CN S0N net35 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX12 CN I2 VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX11 DN I3 VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX10 net44 net35 VSS VPW NHVT11LL_CKT W=0.41u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX5 AN S0N net63 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX7 BN S0 net63 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX8 net48 net63 VSS VPW NHVT11LL_CKT W=0.41u L=40.00n
XX28 S0N S0 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX27 S1N S1 VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX25 ZN net23 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX23 net48 S1 net23 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX21 net44 S1N net23 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX19 DN S0N net35 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX18 CN S0 net35 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX17 CN I2 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX16 DN I3 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX15 net44 net35 VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX9 net48 net63 VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX4 AN S0 net63 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX6 BN S0N net63 VNW PHVT11LL_CKT W=0.5u L=40.00n
.ENDS MUX4NV6_12TH40
.SUBCKT MUX4V0_12TH40 I0 I1 I2 I3 S0 S1 Z VDD VSS
XX7 BN S0 net79 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX5 AN S0N net79 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX11 DN I3 VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX12 CN I2 VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX13 CN S0N net99 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX14 DN S0 net99 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX20 net99 S1 net67 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX22 net79 S1N net67 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX24 Z net67 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX26 S1N S1 VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX29 S0N S0 VSS VPW NHVT11LL_CKT W=0.37u L=40.00n
XX6 BN S0N net79 VNW PHVT11LL_CKT W=0.25u L=40.00n
XX4 AN S0 net79 VNW PHVT11LL_CKT W=0.25u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX16 DN I3 VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX17 CN I2 VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX18 CN S0 net99 VNW PHVT11LL_CKT W=0.25u L=40.00n
XX19 DN S0N net99 VNW PHVT11LL_CKT W=0.25u L=40.00n
XX21 net99 S1N net67 VNW PHVT11LL_CKT W=0.25u L=40.00n
XX23 net79 S1 net67 VNW PHVT11LL_CKT W=0.25u L=40.00n
XX25 Z net67 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX27 S1N S1 VDD VNW PHVT11LL_CKT W=0.24u L=40.00n
XX28 S0N S0 VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
.ENDS MUX4V0_12TH40
.SUBCKT MUX4V1_12TH40 I0 I1 I2 I3 S0 S1 Z VDD VSS
XX7 BN S0 net79 VPW NHVT11LL_CKT W=0.28u L=40.00n
XX5 AN S0N net79 VPW NHVT11LL_CKT W=0.28u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX11 DN I3 VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX12 CN I2 VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX13 CN S0N net99 VPW NHVT11LL_CKT W=0.28u L=40.00n
XX14 DN S0 net99 VPW NHVT11LL_CKT W=0.28u L=40.00n
XX20 net99 S1 net67 VPW NHVT11LL_CKT W=0.28u L=40.00n
XX22 net79 S1N net67 VPW NHVT11LL_CKT W=0.28u L=40.00n
XX24 Z net67 VSS VPW NHVT11LL_CKT W=0.375u L=40.00n
XX26 S1N S1 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX29 S0N S0 VSS VPW NHVT11LL_CKT W=0.46u L=40.00n
XX6 BN S0N net79 VNW PHVT11LL_CKT W=0.35u L=40.00n
XX4 AN S0 net79 VNW PHVT11LL_CKT W=0.35u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX16 DN I3 VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX17 CN I2 VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX18 CN S0 net99 VNW PHVT11LL_CKT W=0.35u L=40.00n
XX19 DN S0N net99 VNW PHVT11LL_CKT W=0.35u L=40.00n
XX21 net99 S1N net67 VNW PHVT11LL_CKT W=0.35u L=40.00n
XX23 net79 S1 net67 VNW PHVT11LL_CKT W=0.35u L=40.00n
XX25 Z net67 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX27 S1N S1 VDD VNW PHVT11LL_CKT W=0.29u L=40.00n
XX28 S0N S0 VDD VNW PHVT11LL_CKT W=0.52u L=40.00n
.ENDS MUX4V1_12TH40
.SUBCKT MUX4V2_12TH40 I0 I1 I2 I3 S0 S1 Z VDD VSS
XX7 BN S0 net79 VPW NHVT11LL_CKT W=335.00n L=40.00n
XX5 AN S0N net79 VPW NHVT11LL_CKT W=335.00n L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=335.00n L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=335.00n L=40.00n
XX11 DN I3 VSS VPW NHVT11LL_CKT W=335.00n L=40.00n
XX12 CN I2 VSS VPW NHVT11LL_CKT W=335.00n L=40.00n
XX13 CN S0N net99 VPW NHVT11LL_CKT W=335.00n L=40.00n
XX14 DN S0 net99 VPW NHVT11LL_CKT W=335.00n L=40.00n
XX20 net99 S1 net67 VPW NHVT11LL_CKT W=335.00n L=40.00n
XX22 net79 S1N net67 VPW NHVT11LL_CKT W=335.00n L=40.00n
XX24 Z net67 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX26 S1N S1 VSS VPW NHVT11LL_CKT W=280.00n L=40.00n
XX29 S0N S0 VSS VPW NHVT11LL_CKT W=520.00n L=40.00n
XX6 BN S0N net79 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX4 AN S0 net79 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX16 DN I3 VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX17 CN I2 VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX18 CN S0 net99 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX19 DN S0N net99 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX21 net99 S1N net67 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX23 net79 S1 net67 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX25 Z net67 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX27 S1N S1 VDD VNW PHVT11LL_CKT W=320.00n L=40.00n
XX28 S0N S0 VDD VNW PHVT11LL_CKT W=590.00n L=40.00n
.ENDS MUX4V2_12TH40
.SUBCKT MUX4V3_12TH40 I0 I1 I2 I3 S0 S1 Z VDD VSS
XX7 BN S0 net79 VPW NHVT11LL_CKT W=0.395u L=40.00n
XX5 AN S0N net79 VPW NHVT11LL_CKT W=0.395u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=0.485u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=0.485u L=40.00n
XX11 DN I3 VSS VPW NHVT11LL_CKT W=0.485u L=40.00n
XX12 CN I2 VSS VPW NHVT11LL_CKT W=0.485u L=40.00n
XX13 CN S0N net99 VPW NHVT11LL_CKT W=0.395u L=40.00n
XX14 DN S0 net99 VPW NHVT11LL_CKT W=0.395u L=40.00n
XX20 net99 S1 net67 VPW NHVT11LL_CKT W=0.395u L=40.00n
XX22 net79 S1N net67 VPW NHVT11LL_CKT W=0.395u L=40.00n
XX24 Z net67 VSS VPW NHVT11LL_CKT W=0.75u L=40.00n
XX26 S1N S1 VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX29 S0N S0 VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX6 BN S0N net79 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX4 AN S0 net79 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX16 DN I3 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX17 CN I2 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX18 CN S0 net99 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX19 DN S0N net99 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX21 net99 S1N net67 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX23 net79 S1 net67 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX25 Z net67 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX27 S1N S1 VDD VNW PHVT11LL_CKT W=0.355u L=40.00n
XX28 S0N S0 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
.ENDS MUX4V3_12TH40
.SUBCKT MUX4V4_12TH40 I0 I1 I2 I3 S0 S1 Z VDD VSS
XX7 BN S0 net79 VPW NHVT11LL_CKT W=0.69u L=40.00n
XX5 AN S0N net79 VPW NHVT11LL_CKT W=0.69u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=0.69u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=0.69u L=40.00n
XX11 DN I3 VSS VPW NHVT11LL_CKT W=0.69u L=40.00n
XX12 CN I2 VSS VPW NHVT11LL_CKT W=0.69u L=40.00n
XX13 CN S0N net99 VPW NHVT11LL_CKT W=0.69u L=40.00n
XX14 DN S0 net99 VPW NHVT11LL_CKT W=0.69u L=40.00n
XX20 net99 S1 net67 VPW NHVT11LL_CKT W=0.69u L=40.00n
XX22 net79 S1N net67 VPW NHVT11LL_CKT W=0.69u L=40.00n
XX24 Z net67 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX26 S1N S1 VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX29 S0N S0 VSS VPW NHVT11LL_CKT W=0.95u L=40.00n
XX6 BN S0N net79 VNW PHVT11LL_CKT W=0.87u L=40.00n
XX4 AN S0 net79 VNW PHVT11LL_CKT W=0.87u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=0.87u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=0.87u L=40.00n
XX16 DN I3 VDD VNW PHVT11LL_CKT W=0.87u L=40.00n
XX17 CN I2 VDD VNW PHVT11LL_CKT W=0.87u L=40.00n
XX18 CN S0 net99 VNW PHVT11LL_CKT W=0.87u L=40.00n
XX19 DN S0N net99 VNW PHVT11LL_CKT W=0.87u L=40.00n
XX21 net99 S1N net67 VNW PHVT11LL_CKT W=0.87u L=40.00n
XX23 net79 S1 net67 VNW PHVT11LL_CKT W=0.87u L=40.00n
XX25 Z net67 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX27 S1N S1 VDD VNW PHVT11LL_CKT W=0.58u L=40.00n
XX28 S0N S0 VDD VNW PHVT11LL_CKT W=1.09u L=40.00n
.ENDS MUX4V4_12TH40
.SUBCKT MUX4V6_12TH40 I0 I1 I2 I3 S0 S1 Z VDD VSS
XX7 BN S0 net79 VPW NHVT11LL_CKT W=0.79u L=40.00n
XX5 AN S0N net79 VPW NHVT11LL_CKT W=0.79u L=40.00n
XX2 AN I0 VSS VPW NHVT11LL_CKT W=0.79u L=40.00n
XX1 BN I1 VSS VPW NHVT11LL_CKT W=0.79u L=40.00n
XX11 DN I3 VSS VPW NHVT11LL_CKT W=0.79u L=40.00n
XX12 CN I2 VSS VPW NHVT11LL_CKT W=0.79u L=40.00n
XX13 CN S0N net99 VPW NHVT11LL_CKT W=0.79u L=40.00n
XX14 DN S0 net99 VPW NHVT11LL_CKT W=0.79u L=40.00n
XX20 net99 S1 net67 VPW NHVT11LL_CKT W=0.79u L=40.00n
XX22 net79 S1N net67 VPW NHVT11LL_CKT W=0.79u L=40.00n
XX24 Z net67 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX26 S1N S1 VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX29 S0N S0 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX6 BN S0N net79 VNW PHVT11LL_CKT W=1u L=40.00n
XX4 AN S0 net79 VNW PHVT11LL_CKT W=1u L=40.00n
XX3 AN I0 VDD VNW PHVT11LL_CKT W=1u L=40.00n
XX0 BN I1 VDD VNW PHVT11LL_CKT W=1u L=40.00n
XX16 DN I3 VDD VNW PHVT11LL_CKT W=1u L=40.00n
XX17 CN I2 VDD VNW PHVT11LL_CKT W=1u L=40.00n
XX18 CN S0 net99 VNW PHVT11LL_CKT W=1u L=40.00n
XX19 DN S0N net99 VNW PHVT11LL_CKT W=1u L=40.00n
XX21 net99 S1N net67 VNW PHVT11LL_CKT W=1u L=40.00n
XX23 net79 S1 net67 VNW PHVT11LL_CKT W=1u L=40.00n
XX25 Z net67 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX27 S1N S1 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX28 S0N S0 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS MUX4V6_12TH40
.SUBCKT NAND2BV0_12TH40 A1 B1 ZN VDD VSS
XX5 net16 B1 VSS VPW NHVT11LL_CKT W=0.305u L=40.00n
XX2 ZN net24 net16 VPW NHVT11LL_CKT W=0.305u L=40.00n
XX0 net24 A1 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX4 ZN B1 VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX3 net24 A1 VDD VNW PHVT11LL_CKT W=0.135u L=40.00n
XX1 ZN net24 VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
.ENDS NAND2BV0_12TH40
.SUBCKT NAND2BV12_12TH40 A1 B1 ZN VDD VSS
XX5 net16 B1 VSS VPW NHVT11LL_CKT W=3.66u L=40.00n
XX2 ZN net24 net16 VPW NHVT11LL_CKT W=3.66u L=40.00n
XX0 net24 A1 VSS VPW NHVT11LL_CKT W=0.8u L=40.00n
XX4 ZN B1 VDD VNW PHVT11LL_CKT W=2.37u L=40.00n
XX3 net24 A1 VDD VNW PHVT11LL_CKT W=0.91u L=40.00n
XX1 ZN net24 VDD VNW PHVT11LL_CKT W=2.37u L=40.00n
.ENDS NAND2BV12_12TH40
.SUBCKT NAND2BV16_12TH40 A1 B1 ZN VDD VSS
XX5 net16 B1 VSS VPW NHVT11LL_CKT W=4.88u L=40.00n
XX2 ZN net24 net16 VPW NHVT11LL_CKT W=4.88u L=40.00n
XX0 net24 A1 VSS VPW NHVT11LL_CKT W=1.05u L=40.00n
XX4 ZN B1 VDD VNW PHVT11LL_CKT W=3.16u L=40.00n
XX3 net24 A1 VDD VNW PHVT11LL_CKT W=1.2u L=40.00n
XX1 ZN net24 VDD VNW PHVT11LL_CKT W=3.16u L=40.00n
.ENDS NAND2BV16_12TH40
.SUBCKT NAND2BV1_12TH40 A1 B1 ZN VDD VSS
XX5 net16 B1 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX2 ZN net24 net16 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX0 net24 A1 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX4 ZN B1 VDD VNW PHVT11LL_CKT W=0.28u L=40.00n
XX3 net24 A1 VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX1 ZN net24 VDD VNW PHVT11LL_CKT W=0.28u L=40.00n
.ENDS NAND2BV1_12TH40
.SUBCKT NAND2BV2_12TH40 A1 B1 ZN VDD VSS
XX5 net16 B1 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX2 ZN net24 net16 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX0 net24 A1 VSS VPW NHVT11LL_CKT W=155.00n L=40.00n
XX4 ZN B1 VDD VNW PHVT11LL_CKT W=395.00n L=40.00n
XX3 net24 A1 VDD VNW PHVT11LL_CKT W=180.00n L=40.00n
XX1 ZN net24 VDD VNW PHVT11LL_CKT W=395.00n L=40.00n
.ENDS NAND2BV2_12TH40
.SUBCKT NAND2BV3_12TH40 A1 B1 ZN VDD VSS
XX5 net16 B1 VSS VPW NHVT11LL_CKT W=0.86u L=40.00n
XX2 ZN net24 net16 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX0 net24 A1 VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX4 ZN B1 VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX3 net24 A1 VDD VNW PHVT11LL_CKT W=0.24u L=40.00n
XX1 ZN net24 VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
.ENDS NAND2BV3_12TH40
.SUBCKT NAND2BV4_12TH40 A1 B1 ZN VDD VSS
XX5 net16 B1 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX2 ZN net24 net16 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX0 net24 A1 VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX4 ZN B1 VDD VNW PHVT11LL_CKT W=0.79u L=40.00n
XX3 net24 A1 VDD VNW PHVT11LL_CKT W=0.32u L=40.00n
XX1 ZN net24 VDD VNW PHVT11LL_CKT W=0.79u L=40.00n
.ENDS NAND2BV4_12TH40
.SUBCKT NAND2BV6_12TH40 A1 B1 ZN VDD VSS
XX5 net16 B1 VSS VPW NHVT11LL_CKT W=1.83u L=40.00n
XX2 ZN net24 net16 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX0 net24 A1 VSS VPW NHVT11LL_CKT W=0.405u L=40.00n
XX4 ZN B1 VDD VNW PHVT11LL_CKT W=1.185u L=40.00n
XX3 net24 A1 VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
XX1 ZN net24 VDD VNW PHVT11LL_CKT W=1.185u L=40.00n
.ENDS NAND2BV6_12TH40
.SUBCKT NAND2BV8_12TH40 A1 B1 ZN VDD VSS
XX5 net16 B1 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX2 ZN net24 net16 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX0 net24 A1 VSS VPW NHVT11LL_CKT W=0.53u L=40.00n
XX4 ZN B1 VDD VNW PHVT11LL_CKT W=1.58u L=40.00n
XX3 net24 A1 VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX1 ZN net24 VDD VNW PHVT11LL_CKT W=1.58u L=40.00n
.ENDS NAND2BV8_12TH40
.SUBCKT NAND2CV0_12TH40 A1 A2 ZN VDD VSS
XX5 net12 A2 VSS VPW NHVT11LL_CKT W=300.00n L=40.00n
XX2 ZN A1 net12 VPW NHVT11LL_CKT W=300.00n L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
XX4 ZN A2 VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
.ENDS NAND2CV0_12TH40
.SUBCKT NAND2CV12_12TH40 A1 A2 ZN VDD VSS
XX5 net12 A2 VSS VPW NHVT11LL_CKT W=3.54u L=40.00n
XX2 ZN A1 net12 VPW NHVT11LL_CKT W=3.54u L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX4 ZN A2 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
.ENDS NAND2CV12_12TH40
.SUBCKT NAND2CV16_12TH40 A1 A2 ZN VDD VSS
XX5 net12 A2 VSS VPW NHVT11LL_CKT W=4.72u L=40.00n
XX2 ZN A1 net12 VPW NHVT11LL_CKT W=4.72u L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX4 ZN A2 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
.ENDS NAND2CV16_12TH40
.SUBCKT NAND2CV1_12TH40 A1 A2 ZN VDD VSS
XX5 net12 A2 VSS VPW NHVT11LL_CKT W=415.00n L=40.00n
XX2 ZN A1 net12 VPW NHVT11LL_CKT W=415.00n L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX4 ZN A2 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
.ENDS NAND2CV1_12TH40
.SUBCKT NAND2CV2_12TH40 A1 A2 ZN VDD VSS
XX5 net12 A2 VSS VPW NHVT11LL_CKT W=590.00n L=40.00n
XX2 ZN A1 net12 VPW NHVT11LL_CKT W=590.00n L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX4 ZN A2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS NAND2CV2_12TH40
.SUBCKT NAND2CV3_12TH40 A1 A2 ZN VDD VSS
XX5 net12 A2 VSS VPW NHVT11LL_CKT W=830.00n L=40.00n
XX2 ZN A1 net12 VPW NHVT11LL_CKT W=830.00n L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX4 ZN A2 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
.ENDS NAND2CV3_12TH40
.SUBCKT NAND2CV4_12TH40 A1 A2 ZN VDD VSS
XX5 net12 A2 VSS VPW NHVT11LL_CKT W=1.18u L=40.00n
XX2 ZN A1 net12 VPW NHVT11LL_CKT W=1.18u L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX4 ZN A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS NAND2CV4_12TH40
.SUBCKT NAND2CV6_12TH40 A1 A2 ZN VDD VSS
XX5 net12 A2 VSS VPW NHVT11LL_CKT W=1.77u L=40.00n
XX2 ZN A1 net12 VPW NHVT11LL_CKT W=1.77u L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX4 ZN A2 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS NAND2CV6_12TH40
.SUBCKT NAND2CV8_12TH40 A1 A2 ZN VDD VSS
XX5 net12 A2 VSS VPW NHVT11LL_CKT W=2.36u L=40.00n
XX2 ZN A1 net12 VPW NHVT11LL_CKT W=2.36u L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX4 ZN A2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS NAND2CV8_12TH40
.SUBCKT NAND2V0_12TH40 A1 A2 ZN VDD VSS
XX5 net12 A2 VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX2 ZN A1 net12 VPW NHVT11LL_CKT W=270.00n L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
XX4 ZN A2 VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
.ENDS NAND2V0_12TH40
.SUBCKT NAND2V12_12TH40 A1 A2 ZN VDD VSS
XX5 net12 A2 VSS VPW NHVT11LL_CKT W=3.24u L=40.00n
XX2 ZN A1 net12 VPW NHVT11LL_CKT W=3.24u L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX4 ZN A2 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
.ENDS NAND2V12_12TH40
.SUBCKT NAND2V16_12TH40 A1 A2 ZN VDD VSS
XX5 net12 A2 VSS VPW NHVT11LL_CKT W=4.32u L=40.00n
XX2 ZN A1 net12 VPW NHVT11LL_CKT W=4.32u L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX4 ZN A2 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
.ENDS NAND2V16_12TH40
.SUBCKT NAND2V1_12TH40 A1 A2 ZN VDD VSS
XX5 net12 A2 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX2 ZN A1 net12 VPW NHVT11LL_CKT W=380.00n L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX4 ZN A2 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
.ENDS NAND2V1_12TH40
.SUBCKT NAND2V2_12TH40 A1 A2 ZN VDD VSS
XX5 net12 A2 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX2 ZN A1 net12 VPW NHVT11LL_CKT W=540.00n L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX4 ZN A2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS NAND2V2_12TH40
.SUBCKT NAND2V3_12TH40 A1 A2 ZN VDD VSS
XX5 net12 A2 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX2 ZN A1 net12 VPW NHVT11LL_CKT W=760.00n L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX4 ZN A2 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
.ENDS NAND2V3_12TH40
.SUBCKT NAND2V4_12TH40 A1 A2 ZN VDD VSS
XX5 net12 A2 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX2 ZN A1 net12 VPW NHVT11LL_CKT W=1.08u L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX4 ZN A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS NAND2V4_12TH40
.SUBCKT NAND2V6_12TH40 A1 A2 ZN VDD VSS
XX5 net12 A2 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX2 ZN A1 net12 VPW NHVT11LL_CKT W=1.62u L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX4 ZN A2 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS NAND2V6_12TH40
.SUBCKT NAND2V8_12TH40 A1 A2 ZN VDD VSS
XX5 net12 A2 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX2 ZN A1 net12 VPW NHVT11LL_CKT W=2.16u L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX4 ZN A2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS NAND2V8_12TH40
.SUBCKT NAND2XBV0_12TH40 A1 B1 ZN VDD VSS
XX0 net12 A1 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX2 ZN B1 net8 VPW NHVT11LL_CKT W=0.305u L=40.00n
XX5 net8 net12 VSS VPW NHVT11LL_CKT W=0.305u L=40.00n
XX3 net12 A1 VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX1 ZN net12 VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX4 ZN B1 VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
.ENDS NAND2XBV0_12TH40
.SUBCKT NAND2XBV12_12TH40 A1 B1 ZN VDD VSS
XX0 net12 A1 VSS VPW NHVT11LL_CKT W=0.8u L=40.00n
XX2 ZN B1 net8 VPW NHVT11LL_CKT W=3.66u L=40.00n
XX5 net8 net12 VSS VPW NHVT11LL_CKT W=3.66u L=40.00n
XX3 net12 A1 VDD VNW PHVT11LL_CKT W=0.91u L=40.00n
XX1 ZN net12 VDD VNW PHVT11LL_CKT W=2.37u L=40.00n
XX4 ZN B1 VDD VNW PHVT11LL_CKT W=2.37u L=40.00n
.ENDS NAND2XBV12_12TH40
.SUBCKT NAND2XBV16_12TH40 A1 B1 ZN VDD VSS
XX0 net12 A1 VSS VPW NHVT11LL_CKT W=1.05u L=40.00n
XX2 ZN B1 net8 VPW NHVT11LL_CKT W=4.88u L=40.00n
XX5 net8 net12 VSS VPW NHVT11LL_CKT W=4.88u L=40.00n
XX3 net12 A1 VDD VNW PHVT11LL_CKT W=1.2u L=40.00n
XX1 ZN net12 VDD VNW PHVT11LL_CKT W=3.16u L=40.00n
XX4 ZN B1 VDD VNW PHVT11LL_CKT W=3.16u L=40.00n
.ENDS NAND2XBV16_12TH40
.SUBCKT NAND2XBV1_12TH40 A1 B1 ZN VDD VSS
XX0 net12 A1 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX2 ZN B1 net8 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX5 net8 net12 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX3 net12 A1 VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX1 ZN net12 VDD VNW PHVT11LL_CKT W=0.28u L=40.00n
XX4 ZN B1 VDD VNW PHVT11LL_CKT W=0.28u L=40.00n
.ENDS NAND2XBV1_12TH40
.SUBCKT NAND2XBV2_12TH40 A1 B1 ZN VDD VSS
XX0 net12 A1 VSS VPW NHVT11LL_CKT W=155.00n L=40.00n
XX2 ZN B1 net8 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX5 net8 net12 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX3 net12 A1 VDD VNW PHVT11LL_CKT W=180.00n L=40.00n
XX1 ZN net12 VDD VNW PHVT11LL_CKT W=395.00n L=40.00n
XX4 ZN B1 VDD VNW PHVT11LL_CKT W=395.00n L=40.00n
.ENDS NAND2XBV2_12TH40
.SUBCKT NAND2XBV3_12TH40 A1 B1 ZN VDD VSS
XX0 net12 A1 VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX2 ZN B1 net8 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX5 net8 net12 VSS VPW NHVT11LL_CKT W=0.86u L=40.00n
XX3 net12 A1 VDD VNW PHVT11LL_CKT W=0.24u L=40.00n
XX1 ZN net12 VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX4 ZN B1 VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
.ENDS NAND2XBV3_12TH40
.SUBCKT NAND2XBV4_12TH40 A1 B1 ZN VDD VSS
XX0 net12 A1 VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX2 ZN B1 net8 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX5 net8 net12 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX3 net12 A1 VDD VNW PHVT11LL_CKT W=0.32u L=40.00n
XX1 ZN net12 VDD VNW PHVT11LL_CKT W=0.79u L=40.00n
XX4 ZN B1 VDD VNW PHVT11LL_CKT W=0.79u L=40.00n
.ENDS NAND2XBV4_12TH40
.SUBCKT NAND2XBV6_12TH40 A1 B1 ZN VDD VSS
XX0 net12 A1 VSS VPW NHVT11LL_CKT W=0.405u L=40.00n
XX2 ZN B1 net8 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX5 net8 net12 VSS VPW NHVT11LL_CKT W=1.83u L=40.00n
XX3 net12 A1 VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
XX1 ZN net12 VDD VNW PHVT11LL_CKT W=1.185u L=40.00n
XX4 ZN B1 VDD VNW PHVT11LL_CKT W=1.185u L=40.00n
.ENDS NAND2XBV6_12TH40
.SUBCKT NAND2XBV8_12TH40 A1 B1 ZN VDD VSS
XX0 net12 A1 VSS VPW NHVT11LL_CKT W=0.53u L=40.00n
XX2 ZN B1 net8 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX5 net8 net12 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX3 net12 A1 VDD VNW PHVT11LL_CKT W=0.605u L=40.00n
XX1 ZN net12 VDD VNW PHVT11LL_CKT W=1.58u L=40.00n
XX4 ZN B1 VDD VNW PHVT11LL_CKT W=1.58u L=40.00n
.ENDS NAND2XBV8_12TH40
.SUBCKT NAND3BBV0_12TH40 A1 A2 B ZN VDD VSS
XX7 ZN net13 net9 VPW NHVT11LL_CKT W=0.305u L=40.00n
XX6 net9 B VSS VPW NHVT11LL_CKT W=0.305u L=40.00n
XX2 net13 A1 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX5 net13 A2 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX3 ZN net13 VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX1 ZN B VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX0 net13 A1 net32 VNW PHVT11LL_CKT W=0.25u L=40.00n
XX4 net32 A2 VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
.ENDS NAND3BBV0_12TH40
.SUBCKT NAND3BBV12_12TH40 A1 A2 B ZN VDD VSS
XX7 ZN net13 net9 VPW NHVT11LL_CKT W=3.66u L=40.00n
XX6 net9 B VSS VPW NHVT11LL_CKT W=3.66u L=40.00n
XX2 net13 A1 VSS VPW NHVT11LL_CKT W=0.855u L=40.00n
XX5 net13 A2 VSS VPW NHVT11LL_CKT W=0.855u L=40.00n
XX3 ZN net13 VDD VNW PHVT11LL_CKT W=2.37u L=40.00n
XX1 ZN B VDD VNW PHVT11LL_CKT W=2.37u L=40.00n
XX0 net13 A1 net32 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX4 net32 A2 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS NAND3BBV12_12TH40
.SUBCKT NAND3BBV16_12TH40 A1 A2 B ZN VDD VSS
XX7 ZN net13 net9 VPW NHVT11LL_CKT W=4.88u L=40.00n
XX6 net9 B VSS VPW NHVT11LL_CKT W=4.88u L=40.00n
XX2 net13 A1 VSS VPW NHVT11LL_CKT W=1.425u L=40.00n
XX5 net13 A2 VSS VPW NHVT11LL_CKT W=1.425u L=40.00n
XX3 ZN net13 VDD VNW PHVT11LL_CKT W=3.16u L=40.00n
XX1 ZN B VDD VNW PHVT11LL_CKT W=3.16u L=40.00n
XX0 net13 A1 net32 VNW PHVT11LL_CKT W=3.05u L=40.00n
XX4 net32 A2 VDD VNW PHVT11LL_CKT W=3.05u L=40.00n
.ENDS NAND3BBV16_12TH40
.SUBCKT NAND3BBV1_12TH40 A1 A2 B ZN VDD VSS
XX7 ZN net13 net9 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX6 net9 B VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX2 net13 A1 VSS VPW NHVT11LL_CKT W=0.145u L=40.00n
XX5 net13 A2 VSS VPW NHVT11LL_CKT W=0.145u L=40.00n
XX3 ZN net13 VDD VNW PHVT11LL_CKT W=0.28u L=40.00n
XX1 ZN B VDD VNW PHVT11LL_CKT W=0.28u L=40.00n
XX0 net13 A1 net32 VNW PHVT11LL_CKT W=0.31u L=40.00n
XX4 net32 A2 VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
.ENDS NAND3BBV1_12TH40
.SUBCKT NAND3BBV2_12TH40 A1 A2 B ZN VDD VSS
XX7 ZN net13 net9 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX6 net9 B VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX2 net13 A1 VSS VPW NHVT11LL_CKT W=185.00n L=40.00n
XX5 net13 A2 VSS VPW NHVT11LL_CKT W=185.00n L=40.00n
XX3 ZN net13 VDD VNW PHVT11LL_CKT W=395.00n L=40.00n
XX1 ZN B VDD VNW PHVT11LL_CKT W=395.00n L=40.00n
XX0 net13 A1 net32 VNW PHVT11LL_CKT W=395.00n L=40.00n
XX4 net32 A2 VDD VNW PHVT11LL_CKT W=395.00n L=40.00n
.ENDS NAND3BBV2_12TH40
.SUBCKT NAND3BBV3_12TH40 A1 A2 B ZN VDD VSS
XX7 ZN net13 net9 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX6 net9 B VSS VPW NHVT11LL_CKT W=0.86u L=40.00n
XX2 net13 A1 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX5 net13 A2 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX3 ZN net13 VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX1 ZN B VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX0 net13 A1 net32 VNW PHVT11LL_CKT W=0.54u L=40.00n
XX4 net32 A2 VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
.ENDS NAND3BBV3_12TH40
.SUBCKT NAND3BBV4_12TH40 A1 A2 B ZN VDD VSS
XX7 ZN net13 net9 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX6 net9 B VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX2 net13 A1 VSS VPW NHVT11LL_CKT W=0.285u L=40.00n
XX5 net13 A2 VSS VPW NHVT11LL_CKT W=0.285u L=40.00n
XX3 ZN net13 VDD VNW PHVT11LL_CKT W=0.79u L=40.00n
XX1 ZN B VDD VNW PHVT11LL_CKT W=0.79u L=40.00n
XX0 net13 A1 net32 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX4 net32 A2 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
.ENDS NAND3BBV4_12TH40
.SUBCKT NAND3BBV6_12TH40 A1 A2 B ZN VDD VSS
XX7 ZN net13 net9 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX6 net9 B VSS VPW NHVT11LL_CKT W=1.83u L=40.00n
XX2 net13 A1 VSS VPW NHVT11LL_CKT W=0.51u L=40.00n
XX5 net13 A2 VSS VPW NHVT11LL_CKT W=0.51u L=40.00n
XX3 ZN net13 VDD VNW PHVT11LL_CKT W=1.185u L=40.00n
XX1 ZN B VDD VNW PHVT11LL_CKT W=1.185u L=40.00n
XX0 net13 A1 net32 VNW PHVT11LL_CKT W=1.09u L=40.00n
XX4 net32 A2 VDD VNW PHVT11LL_CKT W=1.09u L=40.00n
.ENDS NAND3BBV6_12TH40
.SUBCKT NAND3BBV8_12TH40 A1 A2 B ZN VDD VSS
XX7 ZN net13 net9 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX6 net9 B VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX2 net13 A1 VSS VPW NHVT11LL_CKT W=0.57u L=40.00n
XX5 net13 A2 VSS VPW NHVT11LL_CKT W=0.57u L=40.00n
XX3 ZN net13 VDD VNW PHVT11LL_CKT W=1.58u L=40.00n
XX1 ZN B VDD VNW PHVT11LL_CKT W=1.58u L=40.00n
XX0 net13 A1 net32 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX4 net32 A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS NAND3BBV8_12TH40
.SUBCKT NAND3BV0_12TH40 A1 B1 B2 ZN VDD VSS
XX2 net21 A1 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX6 net29 B1 net25 VPW NHVT11LL_CKT W=0.305u L=40.00n
XX7 ZN net21 net29 VPW NHVT11LL_CKT W=0.305u L=40.00n
XX5 net25 B2 VSS VPW NHVT11LL_CKT W=0.305u L=40.00n
XX4 ZN net21 VDD VNW PHVT11LL_CKT W=0.145u L=40.00n
XX0 net21 A1 VDD VNW PHVT11LL_CKT W=0.135u L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=0.145u L=40.00n
XX3 ZN B1 VDD VNW PHVT11LL_CKT W=0.145u L=40.00n
.ENDS NAND3BV0_12TH40
.SUBCKT NAND3BV12_12TH40 A1 B1 B2 ZN VDD VSS
XX2 net21 A1 VSS VPW NHVT11LL_CKT W=0.72u L=40.00n
XX6 net29 B1 net25 VPW NHVT11LL_CKT W=3.66u L=40.00n
XX7 ZN net21 net29 VPW NHVT11LL_CKT W=3.66u L=40.00n
XX5 net25 B2 VSS VPW NHVT11LL_CKT W=3.66u L=40.00n
XX4 ZN net21 VDD VNW PHVT11LL_CKT W=1.71u L=40.00n
XX0 net21 A1 VDD VNW PHVT11LL_CKT W=0.82u L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=1.71u L=40.00n
XX3 ZN B1 VDD VNW PHVT11LL_CKT W=1.71u L=40.00n
.ENDS NAND3BV12_12TH40
.SUBCKT NAND3BV1_12TH40 A1 B1 B2 ZN VDD VSS
XX2 net21 A1 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX6 net29 B1 net25 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX7 ZN net21 net29 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX5 net25 B2 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX4 ZN net21 VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX0 net21 A1 VDD VNW PHVT11LL_CKT W=0.135u L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX3 ZN B1 VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
.ENDS NAND3BV1_12TH40
.SUBCKT NAND3BV2_12TH40 A1 B1 B2 ZN VDD VSS
XX2 net21 A1 VSS VPW NHVT11LL_CKT W=145.00n L=40.00n
XX6 net29 B1 net25 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX7 ZN net21 net29 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX5 net25 B2 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX4 ZN net21 VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX0 net21 A1 VDD VNW PHVT11LL_CKT W=165.00n L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX3 ZN B1 VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
.ENDS NAND3BV2_12TH40
.SUBCKT NAND3BV3_12TH40 A1 B1 B2 ZN VDD VSS
XX2 net21 A1 VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX6 net29 B1 net25 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX7 ZN net21 net29 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX5 net25 B2 VSS VPW NHVT11LL_CKT W=0.86u L=40.00n
XX4 ZN net21 VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX0 net21 A1 VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX3 ZN B1 VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
.ENDS NAND3BV3_12TH40
.SUBCKT NAND3BV4_12TH40 A1 B1 B2 ZN VDD VSS
XX2 net21 A1 VSS VPW NHVT11LL_CKT W=0.255u L=40.00n
XX6 net29 B1 net25 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX7 ZN net21 net29 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX5 net25 B2 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX4 ZN net21 VDD VNW PHVT11LL_CKT W=0.57u L=40.00n
XX0 net21 A1 VDD VNW PHVT11LL_CKT W=0.29u L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=0.57u L=40.00n
XX3 ZN B1 VDD VNW PHVT11LL_CKT W=0.57u L=40.00n
.ENDS NAND3BV4_12TH40
.SUBCKT NAND3BV6_12TH40 A1 B1 B2 ZN VDD VSS
XX2 net21 A1 VSS VPW NHVT11LL_CKT W=0.365u L=40.00n
XX6 net29 B1 net25 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX7 ZN net21 net29 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX5 net25 B2 VSS VPW NHVT11LL_CKT W=1.83u L=40.00n
XX4 ZN net21 VDD VNW PHVT11LL_CKT W=0.855u L=40.00n
XX0 net21 A1 VDD VNW PHVT11LL_CKT W=0.415u L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=0.855u L=40.00n
XX3 ZN B1 VDD VNW PHVT11LL_CKT W=0.855u L=40.00n
.ENDS NAND3BV6_12TH40
.SUBCKT NAND3BV8_12TH40 A1 B1 B2 ZN VDD VSS
XX2 net21 A1 VSS VPW NHVT11LL_CKT W=0.48u L=40.00n
XX6 net29 B1 net25 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX7 ZN net21 net29 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX5 net25 B2 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX4 ZN net21 VDD VNW PHVT11LL_CKT W=1.14u L=40.00n
XX0 net21 A1 VDD VNW PHVT11LL_CKT W=0.545u L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=1.14u L=40.00n
XX3 ZN B1 VDD VNW PHVT11LL_CKT W=1.14u L=40.00n
.ENDS NAND3BV8_12TH40
.SUBCKT NAND3CV0_12TH40 A1 A2 A3 ZN VDD VSS
XX5 net17 A3 VSS VPW NHVT11LL_CKT W=310.00n L=40.00n
XX6 net21 A2 net17 VPW NHVT11LL_CKT W=310.00n L=40.00n
XX7 ZN A1 net21 VPW NHVT11LL_CKT W=310.00n L=40.00n
XX4 ZN A3 VDD VNW PHVT11LL_CKT W=245.00n L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=245.00n L=40.00n
XX3 ZN A2 VDD VNW PHVT11LL_CKT W=245.00n L=40.00n
.ENDS NAND3CV0_12TH40
.SUBCKT NAND3CV12_12TH40 A1 A2 A3 ZN VDD VSS
XX5 net17 A3 VSS VPW NHVT11LL_CKT W=3.66u L=40.00n
XX6 net21 A2 net17 VPW NHVT11LL_CKT W=3.66u L=40.00n
XX7 ZN A1 net21 VPW NHVT11LL_CKT W=3.66u L=40.00n
XX4 ZN A3 VDD VNW PHVT11LL_CKT W=2.88u L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=2.88u L=40.00n
XX3 ZN A2 VDD VNW PHVT11LL_CKT W=2.88u L=40.00n
.ENDS NAND3CV12_12TH40
.SUBCKT NAND3CV1_12TH40 A1 A2 A3 ZN VDD VSS
XX5 net17 A3 VSS VPW NHVT11LL_CKT W=430.00n L=40.00n
XX6 net21 A2 net17 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX7 ZN A1 net21 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX4 ZN A3 VDD VNW PHVT11LL_CKT W=340.00n L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=340.00n L=40.00n
XX3 ZN A2 VDD VNW PHVT11LL_CKT W=340.00n L=40.00n
.ENDS NAND3CV1_12TH40
.SUBCKT NAND3CV2_12TH40 A1 A2 A3 ZN VDD VSS
XX5 net17 A3 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX6 net21 A2 net17 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX7 ZN A1 net21 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX4 ZN A3 VDD VNW PHVT11LL_CKT W=480.00n L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=480.00n L=40.00n
XX3 ZN A2 VDD VNW PHVT11LL_CKT W=480.00n L=40.00n
.ENDS NAND3CV2_12TH40
.SUBCKT NAND3CV3_12TH40 A1 A2 A3 ZN VDD VSS
XX5 net17 A3 VSS VPW NHVT11LL_CKT W=860.00n L=40.00n
XX6 net21 A2 net17 VPW NHVT11LL_CKT W=860.00n L=40.00n
XX7 ZN A1 net21 VPW NHVT11LL_CKT W=860.00n L=40.00n
XX4 ZN A3 VDD VNW PHVT11LL_CKT W=680.00n L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=680.00n L=40.00n
XX3 ZN A2 VDD VNW PHVT11LL_CKT W=680.00n L=40.00n
.ENDS NAND3CV3_12TH40
.SUBCKT NAND3CV4_12TH40 A1 A2 A3 ZN VDD VSS
XX5 net17 A3 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX6 net21 A2 net17 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX7 ZN A1 net21 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX4 ZN A3 VDD VNW PHVT11LL_CKT W=960.00n L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=960.00n L=40.00n
XX3 ZN A2 VDD VNW PHVT11LL_CKT W=960.00n L=40.00n
.ENDS NAND3CV4_12TH40
.SUBCKT NAND3CV6_12TH40 A1 A2 A3 ZN VDD VSS
XX5 net17 A3 VSS VPW NHVT11LL_CKT W=1.83u L=40.00n
XX6 net21 A2 net17 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX7 ZN A1 net21 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX4 ZN A3 VDD VNW PHVT11LL_CKT W=1.44u L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=1.44u L=40.00n
XX3 ZN A2 VDD VNW PHVT11LL_CKT W=1.44u L=40.00n
.ENDS NAND3CV6_12TH40
.SUBCKT NAND3CV8_12TH40 A1 A2 A3 ZN VDD VSS
XX5 net17 A3 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX6 net21 A2 net17 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX7 ZN A1 net21 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX4 ZN A3 VDD VNW PHVT11LL_CKT W=1.92u L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=1.92u L=40.00n
XX3 ZN A2 VDD VNW PHVT11LL_CKT W=1.92u L=40.00n
.ENDS NAND3CV8_12TH40
.SUBCKT NAND3V0_12TH40 A1 A2 A3 ZN VDD VSS
XX7 ZN A1 net9 VPW NHVT11LL_CKT W=270.00n L=40.00n
XX6 net9 A2 net13 VPW NHVT11LL_CKT W=270.00n L=40.00n
XX5 net13 A3 VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX3 ZN A2 VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
XX4 ZN A3 VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
.ENDS NAND3V0_12TH40
.SUBCKT NAND3V12_12TH40 A1 A2 A3 ZN VDD VSS
XX7 ZN A1 net9 VPW NHVT11LL_CKT W=3.24u L=40.00n
XX6 net9 A2 net13 VPW NHVT11LL_CKT W=3.24u L=40.00n
XX5 net13 A3 VSS VPW NHVT11LL_CKT W=3.24u L=40.00n
XX3 ZN A2 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX4 ZN A3 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
.ENDS NAND3V12_12TH40
.SUBCKT NAND3V1_12TH40 A1 A2 A3 ZN VDD VSS
XX7 ZN A1 net9 VPW NHVT11LL_CKT W=380.00n L=40.00n
XX6 net9 A2 net13 VPW NHVT11LL_CKT W=380.00n L=40.00n
XX5 net13 A3 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX3 ZN A2 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX4 ZN A3 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
.ENDS NAND3V1_12TH40
.SUBCKT NAND3V2_12TH40 A1 A2 A3 ZN VDD VSS
XX7 ZN A1 net9 VPW NHVT11LL_CKT W=540.00n L=40.00n
XX6 net9 A2 net13 VPW NHVT11LL_CKT W=540.00n L=40.00n
XX5 net13 A3 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX3 ZN A2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX4 ZN A3 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS NAND3V2_12TH40
.SUBCKT NAND3V3_12TH40 A1 A2 A3 ZN VDD VSS
XX7 ZN A1 net9 VPW NHVT11LL_CKT W=760.00n L=40.00n
XX6 net9 A2 net13 VPW NHVT11LL_CKT W=760.00n L=40.00n
XX5 net13 A3 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX3 ZN A2 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX4 ZN A3 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
.ENDS NAND3V3_12TH40
.SUBCKT NAND3V4_12TH40 A1 A2 A3 ZN VDD VSS
XX7 ZN A1 net9 VPW NHVT11LL_CKT W=1.08u L=40.00n
XX6 net9 A2 net13 VPW NHVT11LL_CKT W=1.08u L=40.00n
XX5 net13 A3 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX3 ZN A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX4 ZN A3 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS NAND3V4_12TH40
.SUBCKT NAND3V6_12TH40 A1 A2 A3 ZN VDD VSS
XX7 ZN A1 net9 VPW NHVT11LL_CKT W=1.62u L=40.00n
XX6 net9 A2 net13 VPW NHVT11LL_CKT W=1.62u L=40.00n
XX5 net13 A3 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX3 ZN A2 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX4 ZN A3 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS NAND3V6_12TH40
.SUBCKT NAND3V8_12TH40 A1 A2 A3 ZN VDD VSS
XX7 ZN A1 net9 VPW NHVT11LL_CKT W=2.16u L=40.00n
XX6 net9 A2 net13 VPW NHVT11LL_CKT W=2.16u L=40.00n
XX5 net13 A3 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX3 ZN A2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 ZN A1 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX4 ZN A3 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS NAND3V8_12TH40
.SUBCKT NAND3XXBV0_12TH40 A1 B1 B2 ZN VDD VSS
XX7 ZN B1 net9 VPW NHVT11LL_CKT W=0.305u L=40.00n
XX6 net9 B2 net13 VPW NHVT11LL_CKT W=0.305u L=40.00n
XX5 net13 net17 VSS VPW NHVT11LL_CKT W=0.305u L=40.00n
XX2 net17 A1 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX3 ZN B2 VDD VNW PHVT11LL_CKT W=0.145u L=40.00n
XX1 ZN B1 VDD VNW PHVT11LL_CKT W=0.145u L=40.00n
XX4 ZN net17 VDD VNW PHVT11LL_CKT W=0.145u L=40.00n
XX0 net17 A1 VDD VNW PHVT11LL_CKT W=0.135u L=40.00n
.ENDS NAND3XXBV0_12TH40
.SUBCKT NAND3XXBV12_12TH40 A1 B1 B2 ZN VDD VSS
XX7 ZN B1 net9 VPW NHVT11LL_CKT W=3.66u L=40.00n
XX6 net9 B2 net13 VPW NHVT11LL_CKT W=3.66u L=40.00n
XX5 net13 net17 VSS VPW NHVT11LL_CKT W=3.66u L=40.00n
XX2 net17 A1 VSS VPW NHVT11LL_CKT W=0.72u L=40.00n
XX3 ZN B2 VDD VNW PHVT11LL_CKT W=1.71u L=40.00n
XX1 ZN B1 VDD VNW PHVT11LL_CKT W=1.71u L=40.00n
XX4 ZN net17 VDD VNW PHVT11LL_CKT W=1.71u L=40.00n
XX0 net17 A1 VDD VNW PHVT11LL_CKT W=0.82u L=40.00n
.ENDS NAND3XXBV12_12TH40
.SUBCKT NAND3XXBV1_12TH40 A1 B1 B2 ZN VDD VSS
XX7 ZN B1 net9 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX6 net9 B2 net13 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX5 net13 net17 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX2 net17 A1 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX3 ZN B2 VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX1 ZN B1 VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX4 ZN net17 VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX0 net17 A1 VDD VNW PHVT11LL_CKT W=0.135u L=40.00n
.ENDS NAND3XXBV1_12TH40
.SUBCKT NAND3XXBV2_12TH40 A1 B1 B2 ZN VDD VSS
XX7 ZN B1 net9 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX6 net9 B2 net13 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX5 net13 net17 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX2 net17 A1 VSS VPW NHVT11LL_CKT W=145.00n L=40.00n
XX3 ZN B2 VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX1 ZN B1 VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX4 ZN net17 VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX0 net17 A1 VDD VNW PHVT11LL_CKT W=165.00n L=40.00n
.ENDS NAND3XXBV2_12TH40
.SUBCKT NAND3XXBV3_12TH40 A1 B1 B2 ZN VDD VSS
XX7 ZN B1 net9 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX6 net9 B2 net13 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX5 net13 net17 VSS VPW NHVT11LL_CKT W=0.86u L=40.00n
XX2 net17 A1 VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX3 ZN B2 VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX1 ZN B1 VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX4 ZN net17 VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX0 net17 A1 VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
.ENDS NAND3XXBV3_12TH40
.SUBCKT NAND3XXBV4_12TH40 A1 B1 B2 ZN VDD VSS
XX7 ZN B1 net9 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX6 net9 B2 net13 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX5 net13 net17 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX2 net17 A1 VSS VPW NHVT11LL_CKT W=0.255u L=40.00n
XX3 ZN B2 VDD VNW PHVT11LL_CKT W=0.57u L=40.00n
XX1 ZN B1 VDD VNW PHVT11LL_CKT W=0.57u L=40.00n
XX4 ZN net17 VDD VNW PHVT11LL_CKT W=0.57u L=40.00n
XX0 net17 A1 VDD VNW PHVT11LL_CKT W=0.29u L=40.00n
.ENDS NAND3XXBV4_12TH40
.SUBCKT NAND3XXBV6_12TH40 A1 B1 B2 ZN VDD VSS
XX7 ZN B1 net9 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX6 net9 B2 net13 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX5 net13 net17 VSS VPW NHVT11LL_CKT W=1.83u L=40.00n
XX2 net17 A1 VSS VPW NHVT11LL_CKT W=0.365u L=40.00n
XX3 ZN B2 VDD VNW PHVT11LL_CKT W=0.855u L=40.00n
XX1 ZN B1 VDD VNW PHVT11LL_CKT W=0.855u L=40.00n
XX4 ZN net17 VDD VNW PHVT11LL_CKT W=0.855u L=40.00n
XX0 net17 A1 VDD VNW PHVT11LL_CKT W=0.415u L=40.00n
.ENDS NAND3XXBV6_12TH40
.SUBCKT NAND3XXBV8_12TH40 A1 B1 B2 ZN VDD VSS
XX7 ZN B1 net9 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX6 net9 B2 net13 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX5 net13 net17 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX2 net17 A1 VSS VPW NHVT11LL_CKT W=0.48u L=40.00n
XX3 ZN B2 VDD VNW PHVT11LL_CKT W=1.14u L=40.00n
XX1 ZN B1 VDD VNW PHVT11LL_CKT W=1.14u L=40.00n
XX4 ZN net17 VDD VNW PHVT11LL_CKT W=1.14u L=40.00n
XX0 net17 A1 VDD VNW PHVT11LL_CKT W=0.545u L=40.00n
.ENDS NAND3XXBV8_12TH40
.SUBCKT NAND4BBV0_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX9 net10 A2 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX8 net10 A1 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX7 ZN net10 net18 VPW NHVT11LL_CKT W=0.305u L=40.00n
XX6 net18 B1 net22 VPW NHVT11LL_CKT W=0.305u L=40.00n
XX5 net22 B2 VSS VPW NHVT11LL_CKT W=0.305u L=40.00n
XX2 net10 A1 net29 VNW PHVT11LL_CKT W=0.26u L=40.00n
XX0 net29 A2 VDD VNW PHVT11LL_CKT W=0.26u L=40.00n
XX3 ZN B1 VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX4 ZN net10 VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
.ENDS NAND4BBV0_12TH40
.SUBCKT NAND4BBV12_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX9 net10 A2 VSS VPW NHVT11LL_CKT W=0.94u L=40.00n
XX8 net10 A1 VSS VPW NHVT11LL_CKT W=0.94u L=40.00n
XX7 ZN net10 net18 VPW NHVT11LL_CKT W=3.66u L=40.00n
XX6 net18 B1 net22 VPW NHVT11LL_CKT W=3.66u L=40.00n
XX5 net22 B2 VSS VPW NHVT11LL_CKT W=3.66u L=40.00n
XX2 net10 A1 net29 VNW PHVT11LL_CKT W=2u L=40.00n
XX0 net29 A2 VDD VNW PHVT11LL_CKT W=2u L=40.00n
XX3 ZN B1 VDD VNW PHVT11LL_CKT W=1.71u L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=1.71u L=40.00n
XX4 ZN net10 VDD VNW PHVT11LL_CKT W=1.71u L=40.00n
.ENDS NAND4BBV12_12TH40
.SUBCKT NAND4BBV1_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX9 net10 A2 VSS VPW NHVT11LL_CKT W=0.135u L=40.00n
XX8 net10 A1 VSS VPW NHVT11LL_CKT W=0.135u L=40.00n
XX7 ZN net10 net18 VPW NHVT11LL_CKT W=0.425u L=40.00n
XX6 net18 B1 net22 VPW NHVT11LL_CKT W=0.425u L=40.00n
XX5 net22 B2 VSS VPW NHVT11LL_CKT W=0.425u L=40.00n
XX2 net10 A1 net29 VNW PHVT11LL_CKT W=0.29u L=40.00n
XX0 net29 A2 VDD VNW PHVT11LL_CKT W=0.29u L=40.00n
XX3 ZN B1 VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX4 ZN net10 VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
.ENDS NAND4BBV1_12TH40
.SUBCKT NAND4BBV2_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX9 net10 A2 VSS VPW NHVT11LL_CKT W=170.00n L=40.00n
XX8 net10 A1 VSS VPW NHVT11LL_CKT W=170.00n L=40.00n
XX7 ZN net10 net18 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX6 net18 B1 net22 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX5 net22 B2 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX2 net10 A1 net29 VNW PHVT11LL_CKT W=365.00n L=40.00n
XX0 net29 A2 VDD VNW PHVT11LL_CKT W=365.00n L=40.00n
XX3 ZN B1 VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX4 ZN net10 VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
.ENDS NAND4BBV2_12TH40
.SUBCKT NAND4BBV3_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX9 net10 A2 VSS VPW NHVT11LL_CKT W=0.225u L=40.00n
XX8 net10 A1 VSS VPW NHVT11LL_CKT W=0.225u L=40.00n
XX7 ZN net10 net18 VPW NHVT11LL_CKT W=0.85u L=40.00n
XX6 net18 B1 net22 VPW NHVT11LL_CKT W=0.85u L=40.00n
XX5 net22 B2 VSS VPW NHVT11LL_CKT W=0.85u L=40.00n
XX2 net10 A1 net29 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX0 net29 A2 VDD VNW PHVT11LL_CKT W=0.48u L=40.00n
XX3 ZN B1 VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX4 ZN net10 VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
.ENDS NAND4BBV3_12TH40
.SUBCKT NAND4BBV4_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX9 net10 A2 VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX8 net10 A1 VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX7 ZN net10 net18 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX6 net18 B1 net22 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX5 net22 B2 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX2 net10 A1 net29 VNW PHVT11LL_CKT W=0.72u L=40.00n
XX0 net29 A2 VDD VNW PHVT11LL_CKT W=0.72u L=40.00n
XX3 ZN B1 VDD VNW PHVT11LL_CKT W=0.57u L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=0.57u L=40.00n
XX4 ZN net10 VDD VNW PHVT11LL_CKT W=0.57u L=40.00n
.ENDS NAND4BBV4_12TH40
.SUBCKT NAND4BBV6_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX9 net10 A2 VSS VPW NHVT11LL_CKT W=0.46u L=40.00n
XX8 net10 A1 VSS VPW NHVT11LL_CKT W=0.46u L=40.00n
XX7 ZN net10 net18 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX6 net18 B1 net22 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX5 net22 B2 VSS VPW NHVT11LL_CKT W=1.83u L=40.00n
XX2 net10 A1 net29 VNW PHVT11LL_CKT W=0.98u L=40.00n
XX0 net29 A2 VDD VNW PHVT11LL_CKT W=0.98u L=40.00n
XX3 ZN B1 VDD VNW PHVT11LL_CKT W=0.855u L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=0.855u L=40.00n
XX4 ZN net10 VDD VNW PHVT11LL_CKT W=0.855u L=40.00n
.ENDS NAND4BBV6_12TH40
.SUBCKT NAND4BBV8_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX9 net10 A2 VSS VPW NHVT11LL_CKT W=0.65u L=40.00n
XX8 net10 A1 VSS VPW NHVT11LL_CKT W=0.65u L=40.00n
XX7 ZN net10 net18 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX6 net18 B1 net22 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX5 net22 B2 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX2 net10 A1 net29 VNW PHVT11LL_CKT W=1.38u L=40.00n
XX0 net29 A2 VDD VNW PHVT11LL_CKT W=1.38u L=40.00n
XX3 ZN B1 VDD VNW PHVT11LL_CKT W=1.14u L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=1.14u L=40.00n
XX4 ZN net10 VDD VNW PHVT11LL_CKT W=1.14u L=40.00n
.ENDS NAND4BBV8_12TH40
.SUBCKT NAND4BV0_12TH40 A1 B1 B2 B3 ZN VDD VSS
XX0 net30 B3 VSS VPW NHVT11LL_CKT W=0.325u L=40.00n
XX5 net34 B2 net30 VPW NHVT11LL_CKT W=0.325u L=40.00n
XX6 net38 B1 net34 VPW NHVT11LL_CKT W=0.325u L=40.00n
XX7 ZN net26 net38 VPW NHVT11LL_CKT W=0.325u L=40.00n
XX8 net26 A1 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX9 ZN B3 VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX4 ZN net26 VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX3 ZN B1 VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX2 net26 A1 VDD VNW PHVT11LL_CKT W=0.135u L=40.00n
.ENDS NAND4BV0_12TH40
.SUBCKT NAND4BV1_12TH40 A1 B1 B2 B3 ZN VDD VSS
XX0 net30 B3 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX5 net34 B2 net30 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX6 net38 B1 net34 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX7 ZN net26 net38 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX8 net26 A1 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX9 ZN B3 VDD VNW PHVT11LL_CKT W=0.16u L=40.00n
XX4 ZN net26 VDD VNW PHVT11LL_CKT W=0.16u L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=0.16u L=40.00n
XX3 ZN B1 VDD VNW PHVT11LL_CKT W=0.16u L=40.00n
XX2 net26 A1 VDD VNW PHVT11LL_CKT W=0.135u L=40.00n
.ENDS NAND4BV1_12TH40
.SUBCKT NAND4BV2_12TH40 A1 B1 B2 B3 ZN VDD VSS
XX0 net30 B3 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX5 net34 B2 net30 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX6 net38 B1 net34 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX7 ZN net26 net38 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX8 net26 A1 VSS VPW NHVT11LL_CKT W=135.00n L=40.00n
XX9 ZN B3 VDD VNW PHVT11LL_CKT W=225.00n L=40.00n
XX4 ZN net26 VDD VNW PHVT11LL_CKT W=225.00n L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=225.00n L=40.00n
XX3 ZN B1 VDD VNW PHVT11LL_CKT W=225.00n L=40.00n
XX2 net26 A1 VDD VNW PHVT11LL_CKT W=155.00n L=40.00n
.ENDS NAND4BV2_12TH40
.SUBCKT NAND4BV3_12TH40 A1 B1 B2 B3 ZN VDD VSS
XX0 net30 B3 VSS VPW NHVT11LL_CKT W=0.86u L=40.00n
XX5 net34 B2 net30 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX6 net38 B1 net34 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX7 ZN net26 net38 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX8 net26 A1 VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX9 ZN B3 VDD VNW PHVT11LL_CKT W=0.32u L=40.00n
XX4 ZN net26 VDD VNW PHVT11LL_CKT W=0.32u L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=0.32u L=40.00n
XX3 ZN B1 VDD VNW PHVT11LL_CKT W=0.32u L=40.00n
XX2 net26 A1 VDD VNW PHVT11LL_CKT W=0.21u L=40.00n
.ENDS NAND4BV3_12TH40
.SUBCKT NAND4BV4_12TH40 A1 B1 B2 B3 ZN VDD VSS
XX0 net30 B3 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX5 net34 B2 net30 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX6 net38 B1 net34 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX7 ZN net26 net38 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX8 net26 A1 VSS VPW NHVT11LL_CKT W=0.24u L=40.00n
XX9 ZN B3 VDD VNW PHVT11LL_CKT W=0.45u L=40.00n
XX4 ZN net26 VDD VNW PHVT11LL_CKT W=0.45u L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=0.45u L=40.00n
XX3 ZN B1 VDD VNW PHVT11LL_CKT W=0.45u L=40.00n
XX2 net26 A1 VDD VNW PHVT11LL_CKT W=0.275u L=40.00n
.ENDS NAND4BV4_12TH40
.SUBCKT NAND4BV6_12TH40 A1 B1 B2 B3 ZN VDD VSS
XX0 net30 B3 VSS VPW NHVT11LL_CKT W=1.83u L=40.00n
XX5 net34 B2 net30 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX6 net38 B1 net34 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX7 ZN net26 net38 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX8 net26 A1 VSS VPW NHVT11LL_CKT W=0.345u L=40.00n
XX9 ZN B3 VDD VNW PHVT11LL_CKT W=0.675u L=40.00n
XX4 ZN net26 VDD VNW PHVT11LL_CKT W=0.675u L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=0.675u L=40.00n
XX3 ZN B1 VDD VNW PHVT11LL_CKT W=0.675u L=40.00n
XX2 net26 A1 VDD VNW PHVT11LL_CKT W=0.39u L=40.00n
.ENDS NAND4BV6_12TH40
.SUBCKT NAND4BV8_12TH40 A1 B1 B2 B3 ZN VDD VSS
XX0 net30 B3 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX5 net34 B2 net30 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX6 net38 B1 net34 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX7 ZN net26 net38 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX8 net26 A1 VSS VPW NHVT11LL_CKT W=0.45u L=40.00n
XX9 ZN B3 VDD VNW PHVT11LL_CKT W=0.9u L=40.00n
XX4 ZN net26 VDD VNW PHVT11LL_CKT W=0.9u L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=0.9u L=40.00n
XX3 ZN B1 VDD VNW PHVT11LL_CKT W=0.9u L=40.00n
XX2 net26 A1 VDD VNW PHVT11LL_CKT W=0.515u L=40.00n
.ENDS NAND4BV8_12TH40
.SUBCKT NAND4CV0_12TH40 A1 A2 A3 A4 ZN VDD VSS
XX7 ZN A1 net10 VPW NHVT11LL_CKT W=310.00n L=40.00n
XX6 net10 A2 net14 VPW NHVT11LL_CKT W=310.00n L=40.00n
XX5 net14 A3 net18 VPW NHVT11LL_CKT W=310.00n L=40.00n
XX0 net18 A4 VSS VPW NHVT11LL_CKT W=310.00n L=40.00n
XX3 ZN A3 VDD VNW PHVT11LL_CKT W=205.00n L=40.00n
XX1 ZN A2 VDD VNW PHVT11LL_CKT W=205.00n L=40.00n
XX4 ZN A4 VDD VNW PHVT11LL_CKT W=205.00n L=40.00n
XX9 ZN A1 VDD VNW PHVT11LL_CKT W=205.00n L=40.00n
.ENDS NAND4CV0_12TH40
.SUBCKT NAND4CV1_12TH40 A1 A2 A3 A4 ZN VDD VSS
XX7 ZN A1 net10 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX6 net10 A2 net14 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX5 net14 A3 net18 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX0 net18 A4 VSS VPW NHVT11LL_CKT W=430.00n L=40.00n
XX3 ZN A3 VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX1 ZN A2 VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX4 ZN A4 VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX9 ZN A1 VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
.ENDS NAND4CV1_12TH40
.SUBCKT NAND4CV2_12TH40 A1 A2 A3 A4 ZN VDD VSS
XX7 ZN A1 net10 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX6 net10 A2 net14 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX5 net14 A3 net18 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX0 net18 A4 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX3 ZN A3 VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX1 ZN A2 VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX4 ZN A4 VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX9 ZN A1 VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
.ENDS NAND4CV2_12TH40
.SUBCKT NAND4CV3_12TH40 A1 A2 A3 A4 ZN VDD VSS
XX7 ZN A1 net10 VPW NHVT11LL_CKT W=860.00n L=40.00n
XX6 net10 A2 net14 VPW NHVT11LL_CKT W=860.00n L=40.00n
XX5 net14 A3 net18 VPW NHVT11LL_CKT W=860.00n L=40.00n
XX0 net18 A4 VSS VPW NHVT11LL_CKT W=860.00n L=40.00n
XX3 ZN A3 VDD VNW PHVT11LL_CKT W=570.00n L=40.00n
XX1 ZN A2 VDD VNW PHVT11LL_CKT W=570.00n L=40.00n
XX4 ZN A4 VDD VNW PHVT11LL_CKT W=570.00n L=40.00n
XX9 ZN A1 VDD VNW PHVT11LL_CKT W=570.00n L=40.00n
.ENDS NAND4CV3_12TH40
.SUBCKT NAND4CV4_12TH40 A1 A2 A3 A4 ZN VDD VSS
XX7 ZN A1 net10 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX6 net10 A2 net14 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX5 net14 A3 net18 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX0 net18 A4 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX3 ZN A3 VDD VNW PHVT11LL_CKT W=800.00n L=40.00n
XX1 ZN A2 VDD VNW PHVT11LL_CKT W=800.00n L=40.00n
XX4 ZN A4 VDD VNW PHVT11LL_CKT W=800.00n L=40.00n
XX9 ZN A1 VDD VNW PHVT11LL_CKT W=800.00n L=40.00n
.ENDS NAND4CV4_12TH40
.SUBCKT NAND4CV6_12TH40 A1 A2 A3 A4 ZN VDD VSS
XX7 ZN A1 net10 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX6 net10 A2 net14 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX5 net14 A3 net18 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX0 net18 A4 VSS VPW NHVT11LL_CKT W=1.83u L=40.00n
XX3 ZN A3 VDD VNW PHVT11LL_CKT W=1.2u L=40.00n
XX1 ZN A2 VDD VNW PHVT11LL_CKT W=1.2u L=40.00n
XX4 ZN A4 VDD VNW PHVT11LL_CKT W=1.2u L=40.00n
XX9 ZN A1 VDD VNW PHVT11LL_CKT W=1.2u L=40.00n
.ENDS NAND4CV6_12TH40
.SUBCKT NAND4CV8_12TH40 A1 A2 A3 A4 ZN VDD VSS
XX7 ZN A1 net10 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX6 net10 A2 net14 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX5 net14 A3 net18 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX0 net18 A4 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX3 ZN A3 VDD VNW PHVT11LL_CKT W=1.6u L=40.00n
XX1 ZN A2 VDD VNW PHVT11LL_CKT W=1.6u L=40.00n
XX4 ZN A4 VDD VNW PHVT11LL_CKT W=1.6u L=40.00n
XX9 ZN A1 VDD VNW PHVT11LL_CKT W=1.6u L=40.00n
.ENDS NAND4CV8_12TH40
.SUBCKT NAND4V0_12TH40 A1 A2 A3 A4 ZN VDD VSS
XX0 net30 A4 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX5 net34 A3 net30 VPW NHVT11LL_CKT W=0.27u L=40.00n
XX6 net38 A2 net34 VPW NHVT11LL_CKT W=0.27u L=40.00n
XX7 ZN A1 net38 VPW NHVT11LL_CKT W=0.27u L=40.00n
XX9 ZN A1 VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX4 ZN A4 VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX1 ZN A2 VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX3 ZN A3 VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
.ENDS NAND4V0_12TH40
.SUBCKT NAND4V1_12TH40 A1 A2 A3 A4 ZN VDD VSS
XX0 net30 A4 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX5 net34 A3 net30 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX6 net38 A2 net34 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX7 ZN A1 net38 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX9 ZN A1 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX4 ZN A4 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX1 ZN A2 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX3 ZN A3 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
.ENDS NAND4V1_12TH40
.SUBCKT NAND4V2_12TH40 A1 A2 A3 A4 ZN VDD VSS
XX0 net30 A4 VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX5 net34 A3 net30 VPW NHVT11LL_CKT W=0.54u L=40.00n
XX6 net38 A2 net34 VPW NHVT11LL_CKT W=0.54u L=40.00n
XX7 ZN A1 net38 VPW NHVT11LL_CKT W=0.54u L=40.00n
XX9 ZN A1 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX4 ZN A4 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX1 ZN A2 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX3 ZN A3 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
.ENDS NAND4V2_12TH40
.SUBCKT NAND4V3_12TH40 A1 A2 A3 A4 ZN VDD VSS
XX0 net30 A4 VSS VPW NHVT11LL_CKT W=0.76u L=40.00n
XX5 net34 A3 net30 VPW NHVT11LL_CKT W=0.76u L=40.00n
XX6 net38 A2 net34 VPW NHVT11LL_CKT W=0.76u L=40.00n
XX7 ZN A1 net38 VPW NHVT11LL_CKT W=0.76u L=40.00n
XX9 ZN A1 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX4 ZN A4 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX1 ZN A2 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX3 ZN A3 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
.ENDS NAND4V3_12TH40
.SUBCKT NAND4V4_12TH40 A1 A2 A3 A4 ZN VDD VSS
XX0 net30 A4 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX5 net34 A3 net30 VPW NHVT11LL_CKT W=1.08u L=40.00n
XX6 net38 A2 net34 VPW NHVT11LL_CKT W=1.08u L=40.00n
XX7 ZN A1 net38 VPW NHVT11LL_CKT W=1.08u L=40.00n
XX9 ZN A1 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX4 ZN A4 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 ZN A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX3 ZN A3 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS NAND4V4_12TH40
.SUBCKT NAND4V6_12TH40 A1 A2 A3 A4 ZN VDD VSS
XX0 net30 A4 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX5 net34 A3 net30 VPW NHVT11LL_CKT W=1.62u L=40.00n
XX6 net38 A2 net34 VPW NHVT11LL_CKT W=1.62u L=40.00n
XX7 ZN A1 net38 VPW NHVT11LL_CKT W=1.62u L=40.00n
XX9 ZN A1 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX4 ZN A4 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX1 ZN A2 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX3 ZN A3 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS NAND4V6_12TH40
.SUBCKT NAND4V8_12TH40 A1 A2 A3 A4 ZN VDD VSS
XX0 net30 A4 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX5 net34 A3 net30 VPW NHVT11LL_CKT W=2.16u L=40.00n
XX6 net38 A2 net34 VPW NHVT11LL_CKT W=2.16u L=40.00n
XX7 ZN A1 net38 VPW NHVT11LL_CKT W=2.16u L=40.00n
XX9 ZN A1 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX4 ZN A4 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 ZN A2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX3 ZN A3 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS NAND4V8_12TH40
.SUBCKT NAND4XXXBV0_12TH40 A1 B1 B2 B3 ZN VDD VSS
XX7 ZN B1 net10 VPW NHVT11LL_CKT W=0.325u L=40.00n
XX6 net10 B2 net14 VPW NHVT11LL_CKT W=0.325u L=40.00n
XX5 net14 B3 net18 VPW NHVT11LL_CKT W=0.325u L=40.00n
XX0 net18 net22 VSS VPW NHVT11LL_CKT W=0.325u L=40.00n
XX8 net22 A1 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX3 ZN B3 VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX4 ZN net22 VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX9 ZN B1 VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX2 net22 A1 VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
.ENDS NAND4XXXBV0_12TH40
.SUBCKT NAND4XXXBV1_12TH40 A1 B1 B2 B3 ZN VDD VSS
XX7 ZN B1 net10 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX6 net10 B2 net14 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX5 net14 B3 net18 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX0 net18 net22 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX8 net22 A1 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX3 ZN B3 VDD VNW PHVT11LL_CKT W=0.16u L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=0.16u L=40.00n
XX4 ZN net22 VDD VNW PHVT11LL_CKT W=0.16u L=40.00n
XX9 ZN B1 VDD VNW PHVT11LL_CKT W=0.16u L=40.00n
XX2 net22 A1 VDD VNW PHVT11LL_CKT W=0.135u L=40.00n
.ENDS NAND4XXXBV1_12TH40
.SUBCKT NAND4XXXBV2_12TH40 A1 B1 B2 B3 ZN VDD VSS
XX7 ZN B1 net10 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX6 net10 B2 net14 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX5 net14 B3 net18 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX0 net18 net22 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX8 net22 A1 VSS VPW NHVT11LL_CKT W=135.00n L=40.00n
XX3 ZN B3 VDD VNW PHVT11LL_CKT W=225.00n L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=225.00n L=40.00n
XX4 ZN net22 VDD VNW PHVT11LL_CKT W=225.00n L=40.00n
XX9 ZN B1 VDD VNW PHVT11LL_CKT W=225.00n L=40.00n
XX2 net22 A1 VDD VNW PHVT11LL_CKT W=155.00n L=40.00n
.ENDS NAND4XXXBV2_12TH40
.SUBCKT NAND4XXXBV3_12TH40 A1 B1 B2 B3 ZN VDD VSS
XX7 ZN B1 net10 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX6 net10 B2 net14 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX5 net14 B3 net18 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX0 net18 net22 VSS VPW NHVT11LL_CKT W=0.86u L=40.00n
XX8 net22 A1 VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX3 ZN B3 VDD VNW PHVT11LL_CKT W=0.32u L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=0.32u L=40.00n
XX4 ZN net22 VDD VNW PHVT11LL_CKT W=0.32u L=40.00n
XX9 ZN B1 VDD VNW PHVT11LL_CKT W=0.32u L=40.00n
XX2 net22 A1 VDD VNW PHVT11LL_CKT W=0.21u L=40.00n
.ENDS NAND4XXXBV3_12TH40
.SUBCKT NAND4XXXBV4_12TH40 A1 B1 B2 B3 ZN VDD VSS
XX7 ZN B1 net10 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX6 net10 B2 net14 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX5 net14 B3 net18 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX0 net18 net22 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX8 net22 A1 VSS VPW NHVT11LL_CKT W=0.24u L=40.00n
XX3 ZN B3 VDD VNW PHVT11LL_CKT W=0.45u L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=0.45u L=40.00n
XX4 ZN net22 VDD VNW PHVT11LL_CKT W=0.45u L=40.00n
XX9 ZN B1 VDD VNW PHVT11LL_CKT W=0.45u L=40.00n
XX2 net22 A1 VDD VNW PHVT11LL_CKT W=0.275u L=40.00n
.ENDS NAND4XXXBV4_12TH40
.SUBCKT NAND4XXXBV6_12TH40 A1 B1 B2 B3 ZN VDD VSS
XX7 ZN B1 net10 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX6 net10 B2 net14 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX5 net14 B3 net18 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX0 net18 net22 VSS VPW NHVT11LL_CKT W=1.83u L=40.00n
XX8 net22 A1 VSS VPW NHVT11LL_CKT W=0.345u L=40.00n
XX3 ZN B3 VDD VNW PHVT11LL_CKT W=0.675u L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=0.675u L=40.00n
XX4 ZN net22 VDD VNW PHVT11LL_CKT W=0.675u L=40.00n
XX9 ZN B1 VDD VNW PHVT11LL_CKT W=0.675u L=40.00n
XX2 net22 A1 VDD VNW PHVT11LL_CKT W=0.39u L=40.00n
.ENDS NAND4XXXBV6_12TH40
.SUBCKT NAND4XXXBV8_12TH40 A1 B1 B2 B3 ZN VDD VSS
XX7 ZN B1 net10 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX6 net10 B2 net14 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX5 net14 B3 net18 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX0 net18 net22 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX8 net22 A1 VSS VPW NHVT11LL_CKT W=0.45u L=40.00n
XX3 ZN B3 VDD VNW PHVT11LL_CKT W=0.9u L=40.00n
XX1 ZN B2 VDD VNW PHVT11LL_CKT W=0.9u L=40.00n
XX4 ZN net22 VDD VNW PHVT11LL_CKT W=0.9u L=40.00n
XX9 ZN B1 VDD VNW PHVT11LL_CKT W=0.9u L=40.00n
XX2 net22 A1 VDD VNW PHVT11LL_CKT W=0.515u L=40.00n
.ENDS NAND4XXXBV8_12TH40
.SUBCKT NDQNV2_12TH40 CKN D QN VDD VSS
XX22 QN net23 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX18 net068 net23 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net23 cn net16 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net16 net068 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net40 c net23 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX9 net32 net40 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net47 c net32 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net40 net47 VSS VPW NHVT11LL_CKT W=360.00n L=40.00n
XX3 net48 cn net47 VPW NHVT11LL_CKT W=150.00n L=40.00n
XX2 net48 D VSS VPW NHVT11LL_CKT W=150.00n L=40.00n
XX23 QN net23 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX21 net068 net23 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net23 c net63 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net63 net068 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net40 cn net23 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=350.00n L=40.00n
XX8 net87 net40 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net47 cn net87 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net40 net47 VDD VNW PHVT11LL_CKT W=0.47u L=40.00n
XX0 net48 c net47 VNW PHVT11LL_CKT W=260.00n L=40.00n
XX1 net48 D VDD VNW PHVT11LL_CKT W=320.00n L=40.00n
.ENDS NDQNV2_12TH40
.SUBCKT NDQNV4_12TH40 CKN D QN VDD VSS
XX22 QN net23 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX18 net068 net23 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net23 cn net16 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net16 net068 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net40 c net23 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX9 net32 net40 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net47 c net32 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net40 net47 VSS VPW NHVT11LL_CKT W=0.39u L=40.00n
XX3 net48 cn net47 VPW NHVT11LL_CKT W=150.00n L=40.00n
XX2 net48 D VSS VPW NHVT11LL_CKT W=150.00n L=40.00n
XX23 QN net23 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX21 net068 net23 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net23 c net63 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net63 net068 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net40 cn net23 VNW PHVT11LL_CKT W=0.44u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=350.00n L=40.00n
XX8 net87 net40 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net47 cn net87 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net40 net47 VDD VNW PHVT11LL_CKT W=0.53u L=40.00n
XX0 net48 c net47 VNW PHVT11LL_CKT W=0.37u L=40.00n
XX1 net48 D VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
.ENDS NDQNV4_12TH40
.SUBCKT NDQNV6_12TH40 CKN D QN VDD VSS
XX22 QN net23 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX18 net068 net23 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net23 cn net16 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net16 net068 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net40 c net23 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX9 net32 net40 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net47 c net32 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net40 net47 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX3 net48 cn net47 VPW NHVT11LL_CKT W=150.00n L=40.00n
XX2 net48 D VSS VPW NHVT11LL_CKT W=150.00n L=40.00n
XX23 QN net23 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX21 net068 net23 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net23 c net63 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net63 net068 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net40 cn net23 VNW PHVT11LL_CKT W=0.52u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=350.00n L=40.00n
XX8 net87 net40 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net47 cn net87 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net40 net47 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net48 c net47 VNW PHVT11LL_CKT W=0.51u L=40.00n
XX1 net48 D VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
.ENDS NDQNV6_12TH40
.SUBCKT NDQV2_12TH40 CKN D Q VDD VSS
XX22 Q net8 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX18 net8 net23 VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX17 net23 cn net16 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net16 net8 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net40 c net23 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX9 net32 net40 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net47 c net32 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net40 net47 VSS VPW NHVT11LL_CKT W=360.00n L=40.00n
XX3 net48 cn net47 VPW NHVT11LL_CKT W=150.00n L=40.00n
XX2 net48 D VSS VPW NHVT11LL_CKT W=150.00n L=40.00n
XX23 Q net8 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX21 net8 net23 VDD VNW PHVT11LL_CKT W=325.00n L=40.00n
XX20 net23 c net63 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net63 net8 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net40 cn net23 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX8 net87 net40 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net47 cn net87 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net40 net47 VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX0 net48 c net47 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX1 net48 D VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
.ENDS NDQV2_12TH40
.SUBCKT NDQV4_12TH40 CKN D Q VDD VSS
XX22 Q net8 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX18 net8 net23 VSS VPW NHVT11LL_CKT W=0.46u L=40.00n
XX17 net23 cn net16 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net16 net8 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net40 c net23 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX9 net32 net40 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net47 c net32 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net40 net47 VSS VPW NHVT11LL_CKT W=0.39u L=40.00n
XX3 net48 cn net47 VPW NHVT11LL_CKT W=150.00n L=40.00n
XX2 net48 D VSS VPW NHVT11LL_CKT W=150.00n L=40.00n
XX23 Q net8 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX21 net8 net23 VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
XX20 net23 c net63 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net63 net8 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net40 cn net23 VNW PHVT11LL_CKT W=0.44u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX8 net87 net40 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net47 cn net87 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net40 net47 VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX0 net48 c net47 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX1 net48 D VDD VNW PHVT11LL_CKT W=0.51u L=40.00n
.ENDS NDQV4_12TH40
.SUBCKT NDQV6_12TH40 CKN D Q VDD VSS
XX22 Q net8 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX18 net8 net23 VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX17 net23 cn net16 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net16 net8 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net40 c net23 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX9 net32 net40 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net47 c net32 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net40 net47 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX3 net48 cn net47 VPW NHVT11LL_CKT W=150.00n L=40.00n
XX2 net48 D VSS VPW NHVT11LL_CKT W=150.00n L=40.00n
XX23 Q net8 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX21 net8 net23 VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX20 net23 c net63 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net63 net8 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net40 cn net23 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX8 net87 net40 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net47 cn net87 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net40 net47 VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX0 net48 c net47 VNW PHVT11LL_CKT W=0.485u L=40.00n
XX1 net48 D VDD VNW PHVT11LL_CKT W=0.565u L=40.00n
.ENDS NDQV6_12TH40
.SUBCKT NDRNQNV2_12TH40 CKN D QN RDN VDD VSS
XX25 net84 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX28 R RDN VSS VPW NHVT11LL_CKT W=210.00n L=40.00n
XX27 net99 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net100 D VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX3 net100 cn net092 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX4 net84 net092 VSS VPW NHVT11LL_CKT W=360.00n L=40.00n
XX6 net092 c net92 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net92 net84 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX14 net84 c net99 VPW NHVT11LL_CKT W=0.26u L=40.00n
XX16 net72 net74 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net99 cn net72 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net74 net99 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net99 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX29 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX26 net19 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX24 net31 R VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX1 net100 D VDD VNW PHVT11LL_CKT W=0.32u L=40.00n
XX0 net100 c net092 VNW PHVT11LL_CKT W=0.26u L=40.00n
XX5 net84 net092 net31 VNW PHVT11LL_CKT W=0.55u L=40.00n
XX7 net092 cn net35 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net35 net84 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX15 net84 cn net99 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX19 net23 net74 net19 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net99 c net23 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net74 net99 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net99 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS NDRNQNV2_12TH40
.SUBCKT NDRNQNV4_12TH40 CKN D QN RDN VDD VSS
XX25 net84 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX28 R RDN VSS VPW NHVT11LL_CKT W=210.00n L=40.00n
XX27 net99 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net100 D VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX3 net100 cn net092 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX4 net84 net092 VSS VPW NHVT11LL_CKT W=0.39u L=40.00n
XX6 net092 c net92 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net92 net84 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX14 net84 c net99 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX16 net72 net74 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net99 cn net72 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net74 net99 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net99 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX29 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX26 net19 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX24 net31 R VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX1 net100 D VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX0 net100 c net092 VNW PHVT11LL_CKT W=0.37u L=40.00n
XX5 net84 net092 net31 VNW PHVT11LL_CKT W=0.55u L=40.00n
XX7 net092 cn net35 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net35 net84 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX15 net84 cn net99 VNW PHVT11LL_CKT W=0.41u L=40.00n
XX19 net23 net74 net19 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net99 c net23 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net74 net99 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net99 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS NDRNQNV4_12TH40
.SUBCKT NDRNQNV6_12TH40 CKN D QN RDN VDD VSS
XX25 net84 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX28 R RDN VSS VPW NHVT11LL_CKT W=210.00n L=40.00n
XX27 net99 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net100 D VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX3 net100 cn net092 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX4 net84 net092 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX6 net092 c net92 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net92 net84 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX14 net84 c net99 VPW NHVT11LL_CKT W=330.00n L=40.00n
XX16 net72 net74 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net99 cn net72 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net74 net99 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net99 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX29 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX26 net19 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX24 net31 R VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX1 net100 D VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net100 c net092 VNW PHVT11LL_CKT W=0.52u L=40.00n
XX5 net84 net092 net31 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX7 net092 cn net35 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net35 net84 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.17u L=40.00n
XX15 net84 cn net99 VNW PHVT11LL_CKT W=0.425u L=40.00n
XX19 net23 net74 net19 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net99 c net23 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net74 net99 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net99 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS NDRNQNV6_12TH40
.SUBCKT NDRNQV2_12TH40 CKN D Q RDN VDD VSS
XX25 net84 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX28 R RDN VSS VPW NHVT11LL_CKT W=210.00n L=40.00n
XX27 net99 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net100 D VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX3 net100 cn net092 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX4 net84 net092 VSS VPW NHVT11LL_CKT W=360.00n L=40.00n
XX6 net092 c net92 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net92 net84 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX14 net84 c net99 VPW NHVT11LL_CKT W=0.26u L=40.00n
XX16 net72 net74 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net99 cn net72 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net74 net99 VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX22 Q net74 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX29 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX26 net19 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX24 net31 R VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX1 net100 D VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX0 net100 c net092 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX5 net84 net092 net31 VNW PHVT11LL_CKT W=0.55u L=40.00n
XX7 net092 cn net35 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net35 net84 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX15 net84 cn net99 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX19 net23 net74 net19 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net99 c net23 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net74 net99 VDD VNW PHVT11LL_CKT W=0.29u L=40.00n
XX23 Q net74 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS NDRNQV2_12TH40
.SUBCKT NDRNQV4_12TH40 CKN D Q RDN VDD VSS
XX25 net84 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX28 R RDN VSS VPW NHVT11LL_CKT W=210.00n L=40.00n
XX27 net99 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net100 D VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX3 net100 cn net092 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX4 net84 net092 VSS VPW NHVT11LL_CKT W=0.39u L=40.00n
XX6 net092 c net92 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net92 net84 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX14 net84 c net99 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX16 net72 net74 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net99 cn net72 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net74 net99 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX22 Q net74 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX29 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX26 net19 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX24 net31 R VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX1 net100 D VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX0 net100 c net092 VNW PHVT11LL_CKT W=0.475u L=40.00n
XX5 net84 net092 net31 VNW PHVT11LL_CKT W=0.55u L=40.00n
XX7 net092 cn net35 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net35 net84 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX15 net84 cn net99 VNW PHVT11LL_CKT W=0.41u L=40.00n
XX19 net23 net74 net19 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net99 c net23 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net74 net99 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX23 Q net74 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS NDRNQV4_12TH40
.SUBCKT NDRNQV6_12TH40 CKN D Q RDN VDD VSS
XX25 net84 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX28 R RDN VSS VPW NHVT11LL_CKT W=210.00n L=40.00n
XX27 net99 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net100 D VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX3 net100 cn net092 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX4 net84 net092 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX6 net092 c net92 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net92 net84 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX14 net84 c net99 VPW NHVT11LL_CKT W=330.00n L=40.00n
XX16 net72 net74 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net99 cn net72 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net74 net99 VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX22 Q net74 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX29 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX26 net19 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX24 net31 R VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX1 net100 D VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net100 c net092 VNW PHVT11LL_CKT W=0.52u L=40.00n
XX5 net84 net092 net31 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX7 net092 cn net35 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net35 net84 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.255u L=40.00n
XX15 net84 cn net99 VNW PHVT11LL_CKT W=0.44u L=40.00n
XX19 net23 net74 net19 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net99 c net23 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net74 net99 VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX23 Q net74 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS NDRNQV6_12TH40
.SUBCKT NDRSNQNV2_12TH40 CKN D QN RDN SDN VDD VSS
XX33 R RDN VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX32 net68 R VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX31 net119 SDN net68 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX29 net76 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX27 net96 R net84 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX26 net84 SDN VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX2 net88 D VSS VPW NHVT11LL_CKT W=150.00n L=40.00n
XX3 net88 cn net0105 VPW NHVT11LL_CKT W=150.00n L=40.00n
XX4 net96 net0105 net84 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX6 net0105 c net104 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net104 net96 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX14 net96 c net119 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX16 net120 net122 net76 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net119 cn net120 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX18 net122 net119 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX22 QN net119 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX34 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX30 net119 SDN VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX28 net55 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX25 net31 R VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX24 net96 SDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX1 net88 D VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX0 net88 c net0105 VNW PHVT11LL_CKT W=0.365u L=40.00n
XX5 net96 net0105 net31 VNW PHVT11LL_CKT W=0.51u L=40.00n
XX7 net0105 cn net35 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net35 net96 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=350.00n L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX15 net96 cn net119 VNW PHVT11LL_CKT W=0.41u L=40.00n
XX19 net59 net122 net55 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net119 c net59 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net122 net119 VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX23 QN net119 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS NDRSNQNV2_12TH40
.SUBCKT NDRSNQNV4_12TH40 CKN D QN RDN SDN VDD VSS
XX33 R RDN VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX32 net68 R VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX31 net119 SDN net68 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX29 net76 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX27 net96 R net84 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX26 net84 SDN VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX2 net88 D VSS VPW NHVT11LL_CKT W=150.00n L=40.00n
XX3 net88 cn net0105 VPW NHVT11LL_CKT W=150.00n L=40.00n
XX4 net96 net0105 net84 VPW NHVT11LL_CKT W=390.00n L=40.00n
XX6 net0105 c net104 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net104 net96 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX14 net96 c net119 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX16 net120 net122 net76 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net119 cn net120 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX18 net122 net119 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX22 QN net119 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX34 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX30 net119 SDN VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX28 net55 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX25 net31 R VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX24 net96 SDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX1 net88 D VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX0 net88 c net0105 VNW PHVT11LL_CKT W=0.485u L=40.00n
XX5 net96 net0105 net31 VNW PHVT11LL_CKT W=0.54u L=40.00n
XX7 net0105 cn net35 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net35 net96 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=350.00n L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX15 net96 cn net119 VNW PHVT11LL_CKT W=0.44u L=40.00n
XX19 net59 net122 net55 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net119 c net59 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net122 net119 VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX23 QN net119 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS NDRSNQNV4_12TH40
.SUBCKT NDRSNQNV6_12TH40 CKN D QN RDN SDN VDD VSS
XX33 R RDN VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX32 net68 R VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX31 net119 SDN net68 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX29 net76 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX27 net96 R net84 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX26 net84 SDN VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX2 net88 D VSS VPW NHVT11LL_CKT W=150.00n L=40.00n
XX3 net88 cn net0105 VPW NHVT11LL_CKT W=150.00n L=40.00n
XX4 net96 net0105 net84 VPW NHVT11LL_CKT W=390.00n L=40.00n
XX6 net0105 c net104 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net104 net96 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX14 net96 c net119 VPW NHVT11LL_CKT W=0.27u L=40.00n
XX16 net120 net122 net76 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net119 cn net120 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX18 net122 net119 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX22 QN net119 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX34 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX30 net119 SDN VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX28 net55 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX25 net31 R VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX24 net96 SDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX1 net88 D VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net88 c net0105 VNW PHVT11LL_CKT W=0.52u L=40.00n
XX5 net96 net0105 net31 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX7 net0105 cn net35 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net35 net96 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=350.00n L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.17u L=40.00n
XX15 net96 cn net119 VNW PHVT11LL_CKT W=0.51u L=40.00n
XX19 net59 net122 net55 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net119 c net59 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net122 net119 VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX23 QN net119 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS NDRSNQNV6_12TH40
.SUBCKT NDRSNQV2_12TH40 CKN D Q RDN SDN VDD VSS
XX33 R RDN VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX32 net68 R VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX31 net119 SDN net68 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX29 net76 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX27 net96 R net84 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX26 net84 SDN VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX2 net88 D VSS VPW NHVT11LL_CKT W=150.00n L=40.00n
XX3 net88 cn net0105 VPW NHVT11LL_CKT W=150.00n L=40.00n
XX4 net96 net0105 net84 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX6 net0105 c net104 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net104 net96 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX14 net96 c net119 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX16 net120 net122 net76 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net119 cn net120 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX18 net122 net119 VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX22 Q net122 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX34 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX30 net119 SDN VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX28 net55 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX25 net31 R VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX24 net96 SDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX1 net88 D VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX0 net88 c net0105 VNW PHVT11LL_CKT W=0.365u L=40.00n
XX5 net96 net0105 net31 VNW PHVT11LL_CKT W=0.51u L=40.00n
XX7 net0105 cn net35 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net35 net96 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX15 net96 cn net119 VNW PHVT11LL_CKT W=0.41u L=40.00n
XX19 net59 net122 net55 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net119 c net59 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net122 net119 VDD VNW PHVT11LL_CKT W=0.29u L=40.00n
XX23 Q net122 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS NDRSNQV2_12TH40
.SUBCKT NDRSNQV4_12TH40 CKN D Q RDN SDN VDD VSS
XX33 R RDN VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX32 net68 R VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX31 net119 SDN net68 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX29 net76 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX27 net96 R net84 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX26 net84 SDN VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX2 net88 D VSS VPW NHVT11LL_CKT W=150.00n L=40.00n
XX3 net88 cn net0105 VPW NHVT11LL_CKT W=150.00n L=40.00n
XX4 net96 net0105 net84 VPW NHVT11LL_CKT W=390.00n L=40.00n
XX6 net0105 c net104 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net104 net96 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX14 net96 c net119 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX16 net120 net122 net76 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net119 cn net120 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX18 net122 net119 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX22 Q net122 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX34 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX30 net119 SDN VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX28 net55 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX25 net31 R VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX24 net96 SDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX1 net88 D VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX0 net88 c net0105 VNW PHVT11LL_CKT W=0.485u L=40.00n
XX5 net96 net0105 net31 VNW PHVT11LL_CKT W=0.54u L=40.00n
XX7 net0105 cn net35 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net35 net96 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX15 net96 cn net119 VNW PHVT11LL_CKT W=0.44u L=40.00n
XX19 net59 net122 net55 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net119 c net59 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net122 net119 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX23 Q net122 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS NDRSNQV4_12TH40
.SUBCKT NDRSNQV6_12TH40 CKN D Q RDN SDN VDD VSS
XX33 R RDN VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX32 net68 R VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX31 net119 SDN net68 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX29 net76 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX27 net96 R net84 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX26 net84 SDN VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX2 net88 D VSS VPW NHVT11LL_CKT W=150.00n L=40.00n
XX3 net88 cn net0105 VPW NHVT11LL_CKT W=150.00n L=40.00n
XX4 net96 net0105 net84 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX6 net0105 c net104 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net104 net96 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX14 net96 c net119 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX16 net120 net122 net76 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net119 cn net120 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX18 net122 net119 VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX22 Q net122 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX34 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX30 net119 SDN VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX28 net55 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX25 net31 R VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX24 net96 SDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX1 net88 D VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net88 c net0105 VNW PHVT11LL_CKT W=0.52u L=40.00n
XX5 net96 net0105 net31 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX7 net0105 cn net35 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net35 net96 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.17u L=40.00n
XX15 net96 cn net119 VNW PHVT11LL_CKT W=0.51u L=40.00n
XX19 net59 net122 net55 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net119 c net59 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net122 net119 VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX23 Q net122 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS NDRSNQV6_12TH40
.SUBCKT NDSNQNV2_12TH40 CKN D QN SDN VDD VSS
XX24 net36 SDN VSS VPW NHVT11LL_CKT W=510.00n L=40.00n
XX22 QN net27 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX18 net14 net27 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net27 cn net12 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX16 net12 net14 net4 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX14 net48 c net27 VPW NHVT11LL_CKT W=0.26u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX9 net28 net48 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net55 c net28 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net48 net55 net36 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX3 net56 cn net55 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX2 net56 D VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX25 net4 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX28 net48 SDN VDD VNW PHVT11LL_CKT W=0.255u L=40.00n
XX29 net27 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net27 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX21 net14 net27 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net27 c net63 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net63 net14 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net48 cn net27 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX8 net91 net48 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net55 cn net91 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net48 net55 VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX0 net56 c net55 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX1 net56 D VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
.ENDS NDSNQNV2_12TH40
.SUBCKT NDSNQNV4_12TH40 CKN D QN SDN VDD VSS
XX24 net36 SDN VSS VPW NHVT11LL_CKT W=510.00n L=40.00n
XX22 QN net27 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX18 net14 net27 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net27 cn net12 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX16 net12 net14 net4 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX14 net48 c net27 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX9 net28 net48 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net55 c net28 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net48 net55 net36 VPW NHVT11LL_CKT W=0.39u L=40.00n
XX3 net56 cn net55 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX2 net56 D VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX25 net4 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX28 net48 SDN VDD VNW PHVT11LL_CKT W=0.225u L=40.00n
XX29 net27 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net27 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX21 net14 net27 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net27 c net63 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net63 net14 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net48 cn net27 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX8 net91 net48 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net55 cn net91 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net48 net55 VDD VNW PHVT11LL_CKT W=0.52u L=40.00n
XX0 net56 c net55 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX1 net56 D VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
.ENDS NDSNQNV4_12TH40
.SUBCKT NDSNQNV6_12TH40 CKN D QN SDN VDD VSS
XX24 net36 SDN VSS VPW NHVT11LL_CKT W=510.00n L=40.00n
XX22 QN net27 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX18 net14 net27 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net27 cn net12 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX16 net12 net14 net4 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX14 net48 c net27 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX9 net28 net48 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net55 c net28 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net48 net55 net36 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX3 net56 cn net55 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX2 net56 D VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX25 net4 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX28 net48 SDN VDD VNW PHVT11LL_CKT W=0.225u L=40.00n
XX29 net27 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net27 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX21 net14 net27 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net27 c net63 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net63 net14 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net48 cn net27 VNW PHVT11LL_CKT W=0.44u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX8 net91 net48 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net55 cn net91 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net48 net55 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net56 c net55 VNW PHVT11LL_CKT W=0.52u L=40.00n
XX1 net56 D VDD VNW PHVT11LL_CKT W=0.59u L=40.00n
.ENDS NDSNQNV6_12TH40
.SUBCKT NDSNQV2_12TH40 CKN D Q SDN VDD VSS
XX24 net36 SDN VSS VPW NHVT11LL_CKT W=510.00n L=40.00n
XX22 Q net14 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX18 net14 net092 VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX17 net092 cn net12 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX16 net12 net14 net4 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX14 net48 c net092 VPW NHVT11LL_CKT W=0.26u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX9 net28 net48 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net55 c net28 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net48 net55 net36 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX3 net56 cn net55 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX2 net56 D VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX25 net4 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX28 net48 SDN VDD VNW PHVT11LL_CKT W=0.225u L=40.00n
XX29 net092 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 Q net14 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX21 net14 net092 VDD VNW PHVT11LL_CKT W=0.29u L=40.00n
XX20 net092 c net63 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net63 net14 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net48 cn net092 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX8 net91 net48 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net55 cn net91 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net48 net55 VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX0 net56 c net55 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX1 net56 D VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
.ENDS NDSNQV2_12TH40
.SUBCKT NDSNQV4_12TH40 CKN D Q SDN VDD VSS
XX24 net36 SDN VSS VPW NHVT11LL_CKT W=510.00n L=40.00n
XX22 Q net14 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX18 net14 net092 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX17 net092 cn net12 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX16 net12 net14 net4 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX14 net48 c net092 VPW NHVT11LL_CKT W=0.39u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX9 net28 net48 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net55 c net28 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net48 net55 net36 VPW NHVT11LL_CKT W=0.39u L=40.00n
XX3 net56 cn net55 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX2 net56 D VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX25 net4 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX28 net48 SDN VDD VNW PHVT11LL_CKT W=0.225u L=40.00n
XX29 net092 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 Q net14 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX21 net14 net092 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX20 net092 c net63 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net63 net14 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net48 cn net092 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX8 net91 net48 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net55 cn net91 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net48 net55 VDD VNW PHVT11LL_CKT W=0.52u L=40.00n
XX0 net56 c net55 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX1 net56 D VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
.ENDS NDSNQV4_12TH40
.SUBCKT NDSNQV6_12TH40 CKN D Q SDN VDD VSS
XX24 net36 SDN VSS VPW NHVT11LL_CKT W=510.00n L=40.00n
XX22 Q net14 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX18 net14 net092 VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX17 net092 cn net12 VPW NHVT11LL_CKT W=0.26u L=40.00n
XX16 net12 net14 net4 VPW NHVT11LL_CKT W=0.26u L=40.00n
XX14 net48 c net092 VPW NHVT11LL_CKT W=330.00n L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX9 net28 net48 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net55 c net28 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net48 net55 net36 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX3 net56 cn net55 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX2 net56 D VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX25 net4 SDN VSS VPW NHVT11LL_CKT W=0.26u L=40.00n
XX28 net48 SDN VDD VNW PHVT11LL_CKT W=0.225u L=40.00n
XX29 net092 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 Q net14 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX21 net14 net092 VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX20 net092 c net63 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net63 net14 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net48 cn net092 VNW PHVT11LL_CKT W=0.455u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX8 net91 net48 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net55 cn net91 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net48 net55 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net56 c net55 VNW PHVT11LL_CKT W=0.52u L=40.00n
XX1 net56 D VDD VNW PHVT11LL_CKT W=0.59u L=40.00n
.ENDS NDSNQV6_12TH40
.SUBCKT NOR2BV0_12TH40 A1 B1 ZN VDD VSS
XX2 ZN B1 VSS VPW NHVT11LL_CKT W=0.145u L=40.00n
XX0 ZN net4 VSS VPW NHVT11LL_CKT W=0.145u L=40.00n
XX4 net4 A1 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX1 ZN net4 net23 VNW PHVT11LL_CKT W=0.305u L=40.00n
XX3 net4 A1 VDD VNW PHVT11LL_CKT W=0.135u L=40.00n
XX9 net23 B1 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
.ENDS NOR2BV0_12TH40
.SUBCKT NOR2BV12_12TH40 A1 B1 ZN VDD VSS
XX2 ZN B1 VSS VPW NHVT11LL_CKT W=1.71u L=40.00n
XX0 ZN net4 VSS VPW NHVT11LL_CKT W=1.71u L=40.00n
XX4 net4 A1 VSS VPW NHVT11LL_CKT W=0.72u L=40.00n
XX1 ZN net4 net23 VNW PHVT11LL_CKT W=3.66u L=40.00n
XX3 net4 A1 VDD VNW PHVT11LL_CKT W=0.82u L=40.00n
XX9 net23 B1 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
.ENDS NOR2BV12_12TH40
.SUBCKT NOR2BV16_12TH40 A1 B1 ZN VDD VSS
XX2 ZN B1 VSS VPW NHVT11LL_CKT W=2.28u L=40.00n
XX0 ZN net4 VSS VPW NHVT11LL_CKT W=2.28u L=40.00n
XX4 net4 A1 VSS VPW NHVT11LL_CKT W=0.95u L=40.00n
XX1 ZN net4 net23 VNW PHVT11LL_CKT W=4.88u L=40.00n
XX3 net4 A1 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX9 net23 B1 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
.ENDS NOR2BV16_12TH40
.SUBCKT NOR2BV1_12TH40 A1 B1 ZN VDD VSS
XX2 ZN B1 VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX0 ZN net4 VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX4 net4 A1 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX1 ZN net4 net23 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX3 net4 A1 VDD VNW PHVT11LL_CKT W=0.135u L=40.00n
XX9 net23 B1 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
.ENDS NOR2BV1_12TH40
.SUBCKT NOR2BV2_12TH40 A1 B1 ZN VDD VSS
XX2 ZN B1 VSS VPW NHVT11LL_CKT W=285.00n L=40.00n
XX0 ZN net4 VSS VPW NHVT11LL_CKT W=285.00n L=40.00n
XX4 net4 A1 VSS VPW NHVT11LL_CKT W=145.00n L=40.00n
XX1 ZN net4 net23 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX3 net4 A1 VDD VNW PHVT11LL_CKT W=165.00n L=40.00n
XX9 net23 B1 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS NOR2BV2_12TH40
.SUBCKT NOR2BV3_12TH40 A1 B1 ZN VDD VSS
XX2 ZN B1 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX0 ZN net4 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX4 net4 A1 VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX1 ZN net4 net23 VNW PHVT11LL_CKT W=0.86u L=40.00n
XX3 net4 A1 VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX9 net23 B1 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
.ENDS NOR2BV3_12TH40
.SUBCKT NOR2BV4_12TH40 A1 B1 ZN VDD VSS
XX2 ZN B1 VSS VPW NHVT11LL_CKT W=0.57u L=40.00n
XX0 ZN net4 VSS VPW NHVT11LL_CKT W=0.57u L=40.00n
XX4 net4 A1 VSS VPW NHVT11LL_CKT W=0.255u L=40.00n
XX1 ZN net4 net23 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX3 net4 A1 VDD VNW PHVT11LL_CKT W=0.29u L=40.00n
XX9 net23 B1 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS NOR2BV4_12TH40
.SUBCKT NOR2BV6_12TH40 A1 B1 ZN VDD VSS
XX2 ZN B1 VSS VPW NHVT11LL_CKT W=0.855u L=40.00n
XX0 ZN net4 VSS VPW NHVT11LL_CKT W=0.855u L=40.00n
XX4 net4 A1 VSS VPW NHVT11LL_CKT W=0.365u L=40.00n
XX1 ZN net4 net23 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX3 net4 A1 VDD VNW PHVT11LL_CKT W=0.415u L=40.00n
XX9 net23 B1 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS NOR2BV6_12TH40
.SUBCKT NOR2BV8_12TH40 A1 B1 ZN VDD VSS
XX2 ZN B1 VSS VPW NHVT11LL_CKT W=1.14u L=40.00n
XX0 ZN net4 VSS VPW NHVT11LL_CKT W=1.14u L=40.00n
XX4 net4 A1 VSS VPW NHVT11LL_CKT W=0.48u L=40.00n
XX1 ZN net4 net23 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX3 net4 A1 VDD VNW PHVT11LL_CKT W=0.545u L=40.00n
XX9 net23 B1 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS NOR2BV8_12TH40
.SUBCKT NOR2CV0_12TH40 A1 A2 ZN VDD VSS
XX2 ZN A1 VSS VPW NHVT11LL_CKT W=140.00n L=40.00n
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=140.00n L=40.00n
XX1 ZN A1 net15 VNW PHVT11LL_CKT W=310.00n L=40.00n
XX9 net15 A2 VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
.ENDS NOR2CV0_12TH40
.SUBCKT NOR2CV12_12TH40 A1 A2 ZN VDD VSS
XX2 ZN A1 VSS VPW NHVT11LL_CKT W=1.65u L=40.00n
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=1.65u L=40.00n
XX1 ZN A1 net15 VNW PHVT11LL_CKT W=3.66u L=40.00n
XX9 net15 A2 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
.ENDS NOR2CV12_12TH40
.SUBCKT NOR2CV16_12TH40 A1 A2 ZN VDD VSS
XX2 ZN A1 VSS VPW NHVT11LL_CKT W=2.2u L=40.00n
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=2.2u L=40.00n
XX1 ZN A1 net15 VNW PHVT11LL_CKT W=4.88u L=40.00n
XX9 net15 A2 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
.ENDS NOR2CV16_12TH40
.SUBCKT NOR2CV1_12TH40 A1 A2 ZN VDD VSS
XX2 ZN A1 VSS VPW NHVT11LL_CKT W=190.00n L=40.00n
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=190.00n L=40.00n
XX1 ZN A1 net15 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX9 net15 A2 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
.ENDS NOR2CV1_12TH40
.SUBCKT NOR2CV2_12TH40 A1 A2 ZN VDD VSS
XX2 ZN A1 VSS VPW NHVT11LL_CKT W=275.00n L=40.00n
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=275.00n L=40.00n
XX1 ZN A1 net15 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX9 net15 A2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS NOR2CV2_12TH40
.SUBCKT NOR2CV3_12TH40 A1 A2 ZN VDD VSS
XX2 ZN A1 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX1 ZN A1 net15 VNW PHVT11LL_CKT W=860.00n L=40.00n
XX9 net15 A2 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
.ENDS NOR2CV3_12TH40
.SUBCKT NOR2CV4_12TH40 A1 A2 ZN VDD VSS
XX2 ZN A1 VSS VPW NHVT11LL_CKT W=550.00n L=40.00n
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=550.00n L=40.00n
XX1 ZN A1 net15 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX9 net15 A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS NOR2CV4_12TH40
.SUBCKT NOR2CV6_12TH40 A1 A2 ZN VDD VSS
XX2 ZN A1 VSS VPW NHVT11LL_CKT W=825.00n L=40.00n
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=825.00n L=40.00n
XX1 ZN A1 net15 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX9 net15 A2 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS NOR2CV6_12TH40
.SUBCKT NOR2CV8_12TH40 A1 A2 ZN VDD VSS
XX2 ZN A1 VSS VPW NHVT11LL_CKT W=1.1u L=40.00n
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=1.1u L=40.00n
XX1 ZN A1 net15 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX9 net15 A2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS NOR2CV8_12TH40
.SUBCKT NOR2V0_12TH40 A1 A2 ZN VDD VSS
XX2 ZN A1 VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX1 ZN A1 net15 VNW PHVT11LL_CKT W=310.00n L=40.00n
XX9 net15 A2 VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
.ENDS NOR2V0_12TH40
.SUBCKT NOR2V12_12TH40 A1 A2 ZN VDD VSS
XX2 ZN A1 VSS VPW NHVT11LL_CKT W=3.24u L=40.00n
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=3.24u L=40.00n
XX1 ZN A1 net15 VNW PHVT11LL_CKT W=3.66u L=40.00n
XX9 net15 A2 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
.ENDS NOR2V12_12TH40
.SUBCKT NOR2V16_12TH40 A1 A2 ZN VDD VSS
XX2 ZN A1 VSS VPW NHVT11LL_CKT W=4.32u L=40.00n
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=4.32u L=40.00n
XX1 ZN A1 net15 VNW PHVT11LL_CKT W=4.88u L=40.00n
XX9 net15 A2 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
.ENDS NOR2V16_12TH40
.SUBCKT NOR2V1_12TH40 A1 A2 ZN VDD VSS
XX2 ZN A1 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX1 ZN A1 net15 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX9 net15 A2 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
.ENDS NOR2V1_12TH40
.SUBCKT NOR2V2_12TH40 A1 A2 ZN VDD VSS
XX2 ZN A1 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX1 ZN A1 net15 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX9 net15 A2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS NOR2V2_12TH40
.SUBCKT NOR2V3_12TH40 A1 A2 ZN VDD VSS
XX2 ZN A1 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX1 ZN A1 net15 VNW PHVT11LL_CKT W=860.00n L=40.00n
XX9 net15 A2 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
.ENDS NOR2V3_12TH40
.SUBCKT NOR2V4_12TH40 A1 A2 ZN VDD VSS
XX2 ZN A1 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX1 ZN A1 net15 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX9 net15 A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS NOR2V4_12TH40
.SUBCKT NOR2V6_12TH40 A1 A2 ZN VDD VSS
XX2 ZN A1 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX1 ZN A1 net15 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX9 net15 A2 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS NOR2V6_12TH40
.SUBCKT NOR2V8_12TH40 A1 A2 ZN VDD VSS
XX2 ZN A1 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX1 ZN A1 net15 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX9 net15 A2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS NOR2V8_12TH40
.SUBCKT NOR2XBV0_12TH40 A1 B1 ZN VDD VSS
XX0 ZN net24 VSS VPW NHVT11LL_CKT W=0.145u L=40.00n
XX2 ZN B1 VSS VPW NHVT11LL_CKT W=0.145u L=40.00n
XX4 net24 A1 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX9 net11 net24 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX1 ZN B1 net11 VNW PHVT11LL_CKT W=0.305u L=40.00n
XX3 net24 A1 VDD VNW PHVT11LL_CKT W=0.135u L=40.00n
.ENDS NOR2XBV0_12TH40
.SUBCKT NOR2XBV12_12TH40 A1 B1 ZN VDD VSS
XX0 ZN net24 VSS VPW NHVT11LL_CKT W=1.71u L=40.00n
XX2 ZN B1 VSS VPW NHVT11LL_CKT W=1.71u L=40.00n
XX4 net24 A1 VSS VPW NHVT11LL_CKT W=0.72u L=40.00n
XX9 net11 net24 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX1 ZN B1 net11 VNW PHVT11LL_CKT W=3.66u L=40.00n
XX3 net24 A1 VDD VNW PHVT11LL_CKT W=0.82u L=40.00n
.ENDS NOR2XBV12_12TH40
.SUBCKT NOR2XBV16_12TH40 A1 B1 ZN VDD VSS
XX0 ZN net24 VSS VPW NHVT11LL_CKT W=2.28u L=40.00n
XX2 ZN B1 VSS VPW NHVT11LL_CKT W=2.28u L=40.00n
XX4 net24 A1 VSS VPW NHVT11LL_CKT W=0.95u L=40.00n
XX9 net11 net24 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX1 ZN B1 net11 VNW PHVT11LL_CKT W=4.88u L=40.00n
XX3 net24 A1 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
.ENDS NOR2XBV16_12TH40
.SUBCKT NOR2XBV1_12TH40 A1 B1 ZN VDD VSS
XX0 ZN net24 VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX2 ZN B1 VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX4 net24 A1 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX9 net11 net24 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX1 ZN B1 net11 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX3 net24 A1 VDD VNW PHVT11LL_CKT W=0.135u L=40.00n
.ENDS NOR2XBV1_12TH40
.SUBCKT NOR2XBV2_12TH40 A1 B1 ZN VDD VSS
XX0 ZN net24 VSS VPW NHVT11LL_CKT W=285.00n L=40.00n
XX2 ZN B1 VSS VPW NHVT11LL_CKT W=285.00n L=40.00n
XX4 net24 A1 VSS VPW NHVT11LL_CKT W=145.00n L=40.00n
XX9 net11 net24 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 ZN B1 net11 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX3 net24 A1 VDD VNW PHVT11LL_CKT W=165.00n L=40.00n
.ENDS NOR2XBV2_12TH40
.SUBCKT NOR2XBV3_12TH40 A1 B1 ZN VDD VSS
XX0 ZN net24 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX2 ZN B1 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX4 net24 A1 VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX9 net11 net24 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX1 ZN B1 net11 VNW PHVT11LL_CKT W=0.86u L=40.00n
XX3 net24 A1 VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
.ENDS NOR2XBV3_12TH40
.SUBCKT NOR2XBV4_12TH40 A1 B1 ZN VDD VSS
XX0 ZN net24 VSS VPW NHVT11LL_CKT W=0.57u L=40.00n
XX2 ZN B1 VSS VPW NHVT11LL_CKT W=0.57u L=40.00n
XX4 net24 A1 VSS VPW NHVT11LL_CKT W=0.255u L=40.00n
XX9 net11 net24 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 ZN B1 net11 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX3 net24 A1 VDD VNW PHVT11LL_CKT W=0.29u L=40.00n
.ENDS NOR2XBV4_12TH40
.SUBCKT NOR2XBV6_12TH40 A1 B1 ZN VDD VSS
XX0 ZN net24 VSS VPW NHVT11LL_CKT W=0.855u L=40.00n
XX2 ZN B1 VSS VPW NHVT11LL_CKT W=0.855u L=40.00n
XX4 net24 A1 VSS VPW NHVT11LL_CKT W=0.365u L=40.00n
XX9 net11 net24 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX1 ZN B1 net11 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX3 net24 A1 VDD VNW PHVT11LL_CKT W=0.415u L=40.00n
.ENDS NOR2XBV6_12TH40
.SUBCKT NOR2XBV8_12TH40 A1 B1 ZN VDD VSS
XX0 ZN net24 VSS VPW NHVT11LL_CKT W=1.14u L=40.00n
XX2 ZN B1 VSS VPW NHVT11LL_CKT W=1.14u L=40.00n
XX4 net24 A1 VSS VPW NHVT11LL_CKT W=0.48u L=40.00n
XX9 net11 net24 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 ZN B1 net11 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX3 net24 A1 VDD VNW PHVT11LL_CKT W=0.545u L=40.00n
.ENDS NOR2XBV8_12TH40
.SUBCKT NOR3BBV0_12TH40 A1 A2 B ZN VDD VSS
XX6 net9 A1 net25 VPW NHVT11LL_CKT W=0.185u L=40.00n
XX4 net25 A2 VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX0 ZN net9 VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX2 ZN B VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX5 net9 A1 VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX3 net9 A2 VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX9 net20 B VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX1 ZN net9 net20 VNW PHVT11LL_CKT W=0.305u L=40.00n
.ENDS NOR3BBV0_12TH40
.SUBCKT NOR3BBV12_12TH40 A1 A2 B ZN VDD VSS
XX6 net9 A1 net25 VPW NHVT11LL_CKT W=1.665u L=40.00n
XX4 net25 A2 VSS VPW NHVT11LL_CKT W=1.665u L=40.00n
XX0 ZN net9 VSS VPW NHVT11LL_CKT W=1.71u L=40.00n
XX2 ZN B VSS VPW NHVT11LL_CKT W=1.71u L=40.00n
XX5 net9 A1 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX3 net9 A2 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX9 net20 B VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX1 ZN net9 net20 VNW PHVT11LL_CKT W=3.66u L=40.00n
.ENDS NOR3BBV12_12TH40
.SUBCKT NOR3BBV16_12TH40 A1 A2 B ZN VDD VSS
XX6 net9 A1 net25 VPW NHVT11LL_CKT W=2.4u L=40.00n
XX4 net25 A2 VSS VPW NHVT11LL_CKT W=2.4u L=40.00n
XX0 ZN net9 VSS VPW NHVT11LL_CKT W=2.28u L=40.00n
XX2 ZN B VSS VPW NHVT11LL_CKT W=2.28u L=40.00n
XX5 net9 A1 VDD VNW PHVT11LL_CKT W=1.56u L=40.00n
XX3 net9 A2 VDD VNW PHVT11LL_CKT W=1.56u L=40.00n
XX9 net20 B VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX1 ZN net9 net20 VNW PHVT11LL_CKT W=4.88u L=40.00n
.ENDS NOR3BBV16_12TH40
.SUBCKT NOR3BBV1_12TH40 A1 A2 B ZN VDD VSS
XX6 net9 A1 net25 VPW NHVT11LL_CKT W=0.235u L=40.00n
XX4 net25 A2 VSS VPW NHVT11LL_CKT W=0.235u L=40.00n
XX0 ZN net9 VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX2 ZN B VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX5 net9 A1 VDD VNW PHVT11LL_CKT W=0.155u L=40.00n
XX3 net9 A2 VDD VNW PHVT11LL_CKT W=0.155u L=40.00n
XX9 net20 B VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX1 ZN net9 net20 VNW PHVT11LL_CKT W=0.425u L=40.00n
.ENDS NOR3BBV1_12TH40
.SUBCKT NOR3BBV2_12TH40 A1 A2 B ZN VDD VSS
XX6 net9 A1 net25 VPW NHVT11LL_CKT W=300.00n L=40.00n
XX4 net25 A2 VSS VPW NHVT11LL_CKT W=300.00n L=40.00n
XX0 ZN net9 VSS VPW NHVT11LL_CKT W=285.00n L=40.00n
XX2 ZN B VSS VPW NHVT11LL_CKT W=285.00n L=40.00n
XX5 net9 A1 VDD VNW PHVT11LL_CKT W=195.00n L=40.00n
XX3 net9 A2 VDD VNW PHVT11LL_CKT W=195.00n L=40.00n
XX9 net20 B VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 ZN net9 net20 VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS NOR3BBV2_12TH40
.SUBCKT NOR3BBV3_12TH40 A1 A2 B ZN VDD VSS
XX6 net9 A1 net25 VPW NHVT11LL_CKT W=0.395u L=40.00n
XX4 net25 A2 VSS VPW NHVT11LL_CKT W=0.395u L=40.00n
XX0 ZN net9 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX2 ZN B VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX5 net9 A1 VDD VNW PHVT11LL_CKT W=0.255u L=40.00n
XX3 net9 A2 VDD VNW PHVT11LL_CKT W=0.255u L=40.00n
XX9 net20 B VDD VNW PHVT11LL_CKT W=0.85u L=40.00n
XX1 ZN net9 net20 VNW PHVT11LL_CKT W=0.85u L=40.00n
.ENDS NOR3BBV3_12TH40
.SUBCKT NOR3BBV4_12TH40 A1 A2 B ZN VDD VSS
XX6 net9 A1 net25 VPW NHVT11LL_CKT W=0.59u L=40.00n
XX4 net25 A2 VSS VPW NHVT11LL_CKT W=0.59u L=40.00n
XX0 ZN net9 VSS VPW NHVT11LL_CKT W=0.57u L=40.00n
XX2 ZN B VSS VPW NHVT11LL_CKT W=0.57u L=40.00n
XX5 net9 A1 VDD VNW PHVT11LL_CKT W=0.385u L=40.00n
XX3 net9 A2 VDD VNW PHVT11LL_CKT W=0.385u L=40.00n
XX9 net20 B VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 ZN net9 net20 VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS NOR3BBV4_12TH40
.SUBCKT NOR3BBV6_12TH40 A1 A2 B ZN VDD VSS
XX6 net9 A1 net25 VPW NHVT11LL_CKT W=0.83u L=40.00n
XX4 net25 A2 VSS VPW NHVT11LL_CKT W=0.83u L=40.00n
XX0 ZN net9 VSS VPW NHVT11LL_CKT W=0.855u L=40.00n
XX2 ZN B VSS VPW NHVT11LL_CKT W=0.855u L=40.00n
XX5 net9 A1 VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX3 net9 A2 VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX9 net20 B VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX1 ZN net9 net20 VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS NOR3BBV6_12TH40
.SUBCKT NOR3BBV8_12TH40 A1 A2 B ZN VDD VSS
XX6 net9 A1 net25 VPW NHVT11LL_CKT W=1.15u L=40.00n
XX4 net25 A2 VSS VPW NHVT11LL_CKT W=1.15u L=40.00n
XX0 ZN net9 VSS VPW NHVT11LL_CKT W=1.14u L=40.00n
XX2 ZN B VSS VPW NHVT11LL_CKT W=1.14u L=40.00n
XX5 net9 A1 VDD VNW PHVT11LL_CKT W=0.75u L=40.00n
XX3 net9 A2 VDD VNW PHVT11LL_CKT W=0.75u L=40.00n
XX9 net20 B VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 ZN net9 net20 VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS NOR3BBV8_12TH40
.SUBCKT NOR3BV1_12TH40 A1 B1 B2 ZN VDD VSS
XX1 net21 A1 VSS VPW NHVT11LL_CKT W=140.00n L=40.00n
XX4 ZN B1 VSS VPW NHVT11LL_CKT W=140.00n L=40.00n
XX5 ZN B2 VSS VPW NHVT11LL_CKT W=140.00n L=40.00n
XX7 ZN net21 VSS VPW NHVT11LL_CKT W=140.00n L=40.00n
XX2 ZN net21 net8 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX3 net8 B1 net12 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX6 net12 B2 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX0 net21 A1 VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
.ENDS NOR3BV1_12TH40
.SUBCKT NOR3BV2_12TH40 A1 B1 B2 ZN VDD VSS
XX1 net21 A1 VSS VPW NHVT11LL_CKT W=200.00n L=40.00n
XX4 ZN B1 VSS VPW NHVT11LL_CKT W=200.00n L=40.00n
XX5 ZN B2 VSS VPW NHVT11LL_CKT W=200.00n L=40.00n
XX7 ZN net21 VSS VPW NHVT11LL_CKT W=200.00n L=40.00n
XX2 ZN net21 net8 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX3 net8 B1 net12 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX6 net12 B2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX0 net21 A1 VDD VNW PHVT11LL_CKT W=230.00n L=40.00n
.ENDS NOR3BV2_12TH40
.SUBCKT NOR3BV4_12TH40 A1 B1 B2 ZN VDD VSS
XX1 net21 A1 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX4 ZN B1 VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX5 ZN B2 VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX7 ZN net21 VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX2 ZN net21 net8 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX3 net8 B1 net12 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX6 net12 B2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 net21 A1 VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
.ENDS NOR3BV4_12TH40
.SUBCKT NOR3BV8_12TH40 A1 B1 B2 ZN VDD VSS
XX1 net21 A1 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX4 ZN B1 VSS VPW NHVT11LL_CKT W=800.00n L=40.00n
XX5 ZN B2 VSS VPW NHVT11LL_CKT W=800.00n L=40.00n
XX7 ZN net21 VSS VPW NHVT11LL_CKT W=800.00n L=40.00n
XX2 ZN net21 net8 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX3 net8 B1 net12 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX6 net12 B2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX0 net21 A1 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS NOR3BV8_12TH40
.SUBCKT NOR3CV0_12TH40 A1 A2 A3 ZN VDD VSS
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 ZN A3 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 ZN A1 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net12 A2 net8 VNW PHVT11LL_CKT W=0.37u L=40.00n
XX1 ZN A1 net12 VNW PHVT11LL_CKT W=0.37u L=40.00n
XX3 net8 A3 VDD VNW PHVT11LL_CKT W=0.37u L=40.00n
.ENDS NOR3CV0_12TH40
.SUBCKT NOR3CV1_12TH40 A1 A2 A3 ZN VDD VSS
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=140.00n L=40.00n
XX2 ZN A3 VSS VPW NHVT11LL_CKT W=140.00n L=40.00n
XX4 ZN A1 VSS VPW NHVT11LL_CKT W=140.00n L=40.00n
XX9 net12 A2 net8 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX1 ZN A1 net12 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX3 net8 A3 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
.ENDS NOR3CV1_12TH40
.SUBCKT NOR3CV2_12TH40 A1 A2 A3 ZN VDD VSS
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=200.00n L=40.00n
XX2 ZN A3 VSS VPW NHVT11LL_CKT W=200.00n L=40.00n
XX4 ZN A1 VSS VPW NHVT11LL_CKT W=200.00n L=40.00n
XX9 net12 A2 net8 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 ZN A1 net12 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX3 net8 A3 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS NOR3CV2_12TH40
.SUBCKT NOR3CV3_12TH40 A1 A2 A3 ZN VDD VSS
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=280.00n L=40.00n
XX2 ZN A3 VSS VPW NHVT11LL_CKT W=280.00n L=40.00n
XX4 ZN A1 VSS VPW NHVT11LL_CKT W=280.00n L=40.00n
XX9 net12 A2 net8 VNW PHVT11LL_CKT W=860.00n L=40.00n
XX1 ZN A1 net12 VNW PHVT11LL_CKT W=860.00n L=40.00n
XX3 net8 A3 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
.ENDS NOR3CV3_12TH40
.SUBCKT NOR3CV4_12TH40 A1 A2 A3 ZN VDD VSS
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX2 ZN A3 VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX4 ZN A1 VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX9 net12 A2 net8 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 ZN A1 net12 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX3 net8 A3 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS NOR3CV4_12TH40
.SUBCKT NOR3CV6_12TH40 A1 A2 A3 ZN VDD VSS
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=600.00n L=40.00n
XX2 ZN A3 VSS VPW NHVT11LL_CKT W=600.00n L=40.00n
XX4 ZN A1 VSS VPW NHVT11LL_CKT W=600.00n L=40.00n
XX9 net12 A2 net8 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX1 ZN A1 net12 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX3 net8 A3 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS NOR3CV6_12TH40
.SUBCKT NOR3CV8_12TH40 A1 A2 A3 ZN VDD VSS
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=800.00n L=40.00n
XX2 ZN A3 VSS VPW NHVT11LL_CKT W=800.00n L=40.00n
XX4 ZN A1 VSS VPW NHVT11LL_CKT W=800.00n L=40.00n
XX9 net12 A2 net8 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 ZN A1 net12 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX3 net8 A3 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS NOR3CV8_12TH40
.SUBCKT NOR3V0_12TH40 A1 A2 A3 ZN VDD VSS
XX4 ZN A1 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX2 ZN A3 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX3 net28 A3 VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX1 ZN A1 net24 VNW PHVT11LL_CKT W=0.31u L=40.00n
XX9 net24 A2 net28 VNW PHVT11LL_CKT W=0.31u L=40.00n
.ENDS NOR3V0_12TH40
.SUBCKT NOR3V1_12TH40 A1 A2 A3 ZN VDD VSS
XX4 ZN A1 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX2 ZN A3 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX3 net28 A3 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX1 ZN A1 net24 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX9 net24 A2 net28 VNW PHVT11LL_CKT W=0.43u L=40.00n
.ENDS NOR3V1_12TH40
.SUBCKT NOR3V2_12TH40 A1 A2 A3 ZN VDD VSS
XX4 ZN A1 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX2 ZN A3 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX3 net28 A3 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 ZN A1 net24 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX9 net24 A2 net28 VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS NOR3V2_12TH40
.SUBCKT NOR3V3_12TH40 A1 A2 A3 ZN VDD VSS
XX4 ZN A1 VSS VPW NHVT11LL_CKT W=0.76u L=40.00n
XX2 ZN A3 VSS VPW NHVT11LL_CKT W=0.76u L=40.00n
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=0.76u L=40.00n
XX3 net28 A3 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX1 ZN A1 net24 VNW PHVT11LL_CKT W=0.86u L=40.00n
XX9 net24 A2 net28 VNW PHVT11LL_CKT W=0.86u L=40.00n
.ENDS NOR3V3_12TH40
.SUBCKT NOR3V4_12TH40 A1 A2 A3 ZN VDD VSS
XX4 ZN A1 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX2 ZN A3 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX3 net28 A3 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 ZN A1 net24 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX9 net24 A2 net28 VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS NOR3V4_12TH40
.SUBCKT NOR3V6_12TH40 A1 A2 A3 ZN VDD VSS
XX4 ZN A1 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX2 ZN A3 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX3 net28 A3 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX1 ZN A1 net24 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX9 net24 A2 net28 VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS NOR3V6_12TH40
.SUBCKT NOR3V8_12TH40 A1 A2 A3 ZN VDD VSS
XX4 ZN A1 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX2 ZN A3 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX0 ZN A2 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX3 net28 A3 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 ZN A1 net24 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX9 net24 A2 net28 VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS NOR3V8_12TH40
.SUBCKT NOR4BBV0_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX8 net26 A2 VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX6 net10 A1 net26 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX0 ZN B1 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX2 ZN B2 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX4 ZN net10 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX7 net10 A1 VDD VNW PHVT11LL_CKT W=0.13u L=40.00n
XX5 net10 A2 VDD VNW PHVT11LL_CKT W=0.13u L=40.00n
XX9 net21 B1 net17 VNW PHVT11LL_CKT W=0.37u L=40.00n
XX1 ZN net10 net21 VNW PHVT11LL_CKT W=0.37u L=40.00n
XX3 net17 B2 VDD VNW PHVT11LL_CKT W=0.37u L=40.00n
.ENDS NOR4BBV0_12TH40
.SUBCKT NOR4BBV1_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX8 net26 A2 VSS VPW NHVT11LL_CKT W=0.225u L=40.00n
XX6 net10 A1 net26 VPW NHVT11LL_CKT W=0.225u L=40.00n
XX0 ZN B1 VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX2 ZN B2 VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX4 ZN net10 VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX7 net10 A1 VDD VNW PHVT11LL_CKT W=0.145u L=40.00n
XX5 net10 A2 VDD VNW PHVT11LL_CKT W=0.145u L=40.00n
XX9 net21 B1 net17 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX1 ZN net10 net21 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX3 net17 B2 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
.ENDS NOR4BBV1_12TH40
.SUBCKT NOR4BBV2_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX8 net26 A2 VSS VPW NHVT11LL_CKT W=280.00n L=40.00n
XX6 net10 A1 net26 VPW NHVT11LL_CKT W=280.00n L=40.00n
XX0 ZN B1 VSS VPW NHVT11LL_CKT W=200.00n L=40.00n
XX2 ZN B2 VSS VPW NHVT11LL_CKT W=200.00n L=40.00n
XX4 ZN net10 VSS VPW NHVT11LL_CKT W=200.00n L=40.00n
XX7 net10 A1 VDD VNW PHVT11LL_CKT W=180.00n L=40.00n
XX5 net10 A2 VDD VNW PHVT11LL_CKT W=180.00n L=40.00n
XX9 net21 B1 net17 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 ZN net10 net21 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX3 net17 B2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS NOR4BBV2_12TH40
.SUBCKT NOR4BBV3_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX8 net26 A2 VSS VPW NHVT11LL_CKT W=0.39u L=40.00n
XX6 net10 A1 net26 VPW NHVT11LL_CKT W=0.39u L=40.00n
XX0 ZN B1 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX2 ZN B2 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX4 ZN net10 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX7 net10 A1 VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX5 net10 A2 VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX9 net21 B1 net17 VNW PHVT11LL_CKT W=0.85u L=40.00n
XX1 ZN net10 net21 VNW PHVT11LL_CKT W=0.85u L=40.00n
XX3 net17 B2 VDD VNW PHVT11LL_CKT W=0.85u L=40.00n
.ENDS NOR4BBV3_12TH40
.SUBCKT NOR4BBV4_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX8 net26 A2 VSS VPW NHVT11LL_CKT W=0.55u L=40.00n
XX6 net10 A1 net26 VPW NHVT11LL_CKT W=0.55u L=40.00n
XX0 ZN B1 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX2 ZN B2 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX4 ZN net10 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX7 net10 A1 VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX5 net10 A2 VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX9 net21 B1 net17 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 ZN net10 net21 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX3 net17 B2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS NOR4BBV4_12TH40
.SUBCKT NOR4BBV6_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX8 net26 A2 VSS VPW NHVT11LL_CKT W=0.77u L=40.00n
XX6 net10 A1 net26 VPW NHVT11LL_CKT W=0.77u L=40.00n
XX0 ZN B1 VSS VPW NHVT11LL_CKT W=0.6u L=40.00n
XX2 ZN B2 VSS VPW NHVT11LL_CKT W=0.6u L=40.00n
XX4 ZN net10 VSS VPW NHVT11LL_CKT W=0.6u L=40.00n
XX7 net10 A1 VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX5 net10 A2 VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX9 net21 B1 net17 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX1 ZN net10 net21 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX3 net17 B2 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS NOR4BBV6_12TH40
.SUBCKT NOR4BBV8_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX8 net26 A2 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX6 net10 A1 net26 VPW NHVT11LL_CKT W=1.07u L=40.00n
XX0 ZN B1 VSS VPW NHVT11LL_CKT W=0.8u L=40.00n
XX2 ZN B2 VSS VPW NHVT11LL_CKT W=0.8u L=40.00n
XX4 ZN net10 VSS VPW NHVT11LL_CKT W=0.8u L=40.00n
XX7 net10 A1 VDD VNW PHVT11LL_CKT W=0.7u L=40.00n
XX5 net10 A2 VDD VNW PHVT11LL_CKT W=0.7u L=40.00n
XX9 net21 B1 net17 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 ZN net10 net21 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX3 net17 B2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS NOR4BBV8_12TH40
.SUBCKT NOR4BV1_12TH40 A1 B1 B2 B3 ZN VDD VSS
XX1 net6 A1 VSS VPW NHVT11LL_CKT W=130.00n L=40.00n
XX7 ZN net6 VSS VPW NHVT11LL_CKT W=130.00n L=40.00n
XX5 ZN B3 VSS VPW NHVT11LL_CKT W=130.00n L=40.00n
XX4 ZN B2 VSS VPW NHVT11LL_CKT W=130.00n L=40.00n
XX8 ZN B1 VSS VPW NHVT11LL_CKT W=130.00n L=40.00n
XX0 net6 A1 VDD VNW PHVT11LL_CKT W=145.00n L=40.00n
XX6 net37 B2 net33 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX3 net41 B1 net37 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX2 ZN net6 net41 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX9 net33 B3 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
.ENDS NOR4BV1_12TH40
.SUBCKT NOR4BV2_12TH40 A1 B1 B2 B3 ZN VDD VSS
XX1 net6 A1 VSS VPW NHVT11LL_CKT W=165.00n L=40.00n
XX7 ZN net6 VSS VPW NHVT11LL_CKT W=165.00n L=40.00n
XX5 ZN B3 VSS VPW NHVT11LL_CKT W=165.00n L=40.00n
XX4 ZN B2 VSS VPW NHVT11LL_CKT W=165.00n L=40.00n
XX8 ZN B1 VSS VPW NHVT11LL_CKT W=165.00n L=40.00n
XX0 net6 A1 VDD VNW PHVT11LL_CKT W=185.00n L=40.00n
XX6 net37 B2 net33 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX3 net41 B1 net37 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX2 ZN net6 net41 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX9 net33 B3 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS NOR4BV2_12TH40
.SUBCKT NOR4BV4_12TH40 A1 B1 B2 B3 ZN VDD VSS
XX1 net6 A1 VSS VPW NHVT11LL_CKT W=330.00n L=40.00n
XX7 ZN net6 VSS VPW NHVT11LL_CKT W=330.00n L=40.00n
XX5 ZN B3 VSS VPW NHVT11LL_CKT W=330.00n L=40.00n
XX4 ZN B2 VSS VPW NHVT11LL_CKT W=330.00n L=40.00n
XX8 ZN B1 VSS VPW NHVT11LL_CKT W=330.00n L=40.00n
XX0 net6 A1 VDD VNW PHVT11LL_CKT W=390.00n L=40.00n
XX6 net37 B2 net33 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX3 net41 B1 net37 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX2 ZN net6 net41 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX9 net33 B3 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS NOR4BV4_12TH40
.SUBCKT NOR4BV8_12TH40 A1 B1 B2 B3 ZN VDD VSS
XX1 net6 A1 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX7 ZN net6 VSS VPW NHVT11LL_CKT W=660.00n L=40.00n
XX5 ZN B3 VSS VPW NHVT11LL_CKT W=660.00n L=40.00n
XX4 ZN B2 VSS VPW NHVT11LL_CKT W=660.00n L=40.00n
XX8 ZN B1 VSS VPW NHVT11LL_CKT W=660.00n L=40.00n
XX0 net6 A1 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX6 net37 B2 net33 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX3 net41 B1 net37 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX2 ZN net6 net41 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX9 net33 B3 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS NOR4BV8_12TH40
.SUBCKT NOR4CV1_12TH40 A1 A2 A3 A4 ZN VDD VSS
XX7 ZN A1 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX5 ZN A4 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 ZN A3 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX8 ZN A2 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net29 A3 net25 VNW PHVT11LL_CKT W=460.00n L=40.00n
XX3 net33 A2 net29 VNW PHVT11LL_CKT W=460.00n L=40.00n
XX2 ZN A1 net33 VNW PHVT11LL_CKT W=460.00n L=40.00n
XX9 net25 A4 VDD VNW PHVT11LL_CKT W=460.00n L=40.00n
.ENDS NOR4CV1_12TH40
.SUBCKT NOR4CV2_12TH40 A1 A2 A3 A4 ZN VDD VSS
XX7 ZN A1 VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX5 ZN A4 VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX4 ZN A3 VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX8 ZN A2 VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX6 net29 A3 net25 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX3 net33 A2 net29 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX2 ZN A1 net33 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX9 net25 A4 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS NOR4CV2_12TH40
.SUBCKT NOR4CV4_12TH40 A1 A2 A3 A4 ZN VDD VSS
XX7 ZN A1 VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX5 ZN A4 VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX4 ZN A3 VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX8 ZN A2 VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX6 net29 A3 net25 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX3 net33 A2 net29 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX2 ZN A1 net33 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX9 net25 A4 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS NOR4CV4_12TH40
.SUBCKT NOR4V1_12TH40 A1 A2 A3 A4 ZN VDD VSS
XX7 ZN A1 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX5 ZN A4 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX4 ZN A3 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX8 ZN A2 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX6 net29 A3 net25 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX3 net33 A2 net29 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX2 ZN A1 net33 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX9 net25 A4 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
.ENDS NOR4V1_12TH40
.SUBCKT NOR4V2_12TH40 A1 A2 A3 A4 ZN VDD VSS
XX7 ZN A1 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX5 ZN A4 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX4 ZN A3 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX8 ZN A2 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX6 net29 A3 net25 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX3 net33 A2 net29 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX2 ZN A1 net33 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX9 net25 A4 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS NOR4V2_12TH40
.SUBCKT NOR4V4_12TH40 A1 A2 A3 A4 ZN VDD VSS
XX7 ZN A1 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX5 ZN A4 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX4 ZN A3 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX8 ZN A2 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX6 net29 A3 net25 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX3 net33 A2 net29 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX2 ZN A1 net33 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX9 net25 A4 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS NOR4V4_12TH40
.SUBCKT OA1B2V0_12TH40 A1 A2 B Z VDD VSS
XX4 net5 A2 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX1 net5 A1 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX2 Z B VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX0 Z net5 VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX5 net24 A2 VDD VNW PHVT11LL_CKT W=0.255u L=40.00n
XX6 net5 A1 net24 VNW PHVT11LL_CKT W=0.255u L=40.00n
XX3 net36 B VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX9 Z net5 net36 VNW PHVT11LL_CKT W=0.305u L=40.00n
.ENDS OA1B2V0_12TH40
.SUBCKT OA1B2V12_12TH40 A1 A2 B Z VDD VSS
XX4 net5 A2 VSS VPW NHVT11LL_CKT W=0.855u L=40.00n
XX1 net5 A1 VSS VPW NHVT11LL_CKT W=0.855u L=40.00n
XX2 Z B VSS VPW NHVT11LL_CKT W=1.71u L=40.00n
XX0 Z net5 VSS VPW NHVT11LL_CKT W=1.71u L=40.00n
XX5 net24 A2 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX6 net5 A1 net24 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX3 net36 B VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX9 Z net5 net36 VNW PHVT11LL_CKT W=3.66u L=40.00n
.ENDS OA1B2V12_12TH40
.SUBCKT OA1B2V16_12TH40 A1 A2 B Z VDD VSS
XX4 net5 A2 VSS VPW NHVT11LL_CKT W=1.35u L=40.00n
XX1 net5 A1 VSS VPW NHVT11LL_CKT W=1.35u L=40.00n
XX2 Z B VSS VPW NHVT11LL_CKT W=2.28u L=40.00n
XX0 Z net5 VSS VPW NHVT11LL_CKT W=2.28u L=40.00n
XX5 net24 A2 VDD VNW PHVT11LL_CKT W=2.9u L=40.00n
XX6 net5 A1 net24 VNW PHVT11LL_CKT W=2.9u L=40.00n
XX3 net36 B VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX9 Z net5 net36 VNW PHVT11LL_CKT W=4.88u L=40.00n
.ENDS OA1B2V16_12TH40
.SUBCKT OA1B2V1_12TH40 A1 A2 B Z VDD VSS
XX4 net5 A2 VSS VPW NHVT11LL_CKT W=0.135u L=40.00n
XX1 net5 A1 VSS VPW NHVT11LL_CKT W=0.135u L=40.00n
XX2 Z B VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX0 Z net5 VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX5 net24 A2 VDD VNW PHVT11LL_CKT W=0.29u L=40.00n
XX6 net5 A1 net24 VNW PHVT11LL_CKT W=0.29u L=40.00n
XX3 net36 B VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX9 Z net5 net36 VNW PHVT11LL_CKT W=0.43u L=40.00n
.ENDS OA1B2V1_12TH40
.SUBCKT OA1B2V2_12TH40 A1 A2 B Z VDD VSS
XX4 net5 A2 VSS VPW NHVT11LL_CKT W=170.00n L=40.00n
XX1 net5 A1 VSS VPW NHVT11LL_CKT W=170.00n L=40.00n
XX2 Z B VSS VPW NHVT11LL_CKT W=285.00n L=40.00n
XX0 Z net5 VSS VPW NHVT11LL_CKT W=285.00n L=40.00n
XX5 net24 A2 VDD VNW PHVT11LL_CKT W=365.00n L=40.00n
XX6 net5 A1 net24 VNW PHVT11LL_CKT W=365.00n L=40.00n
XX3 net36 B VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX9 Z net5 net36 VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS OA1B2V2_12TH40
.SUBCKT OA1B2V3_12TH40 A1 A2 B Z VDD VSS
XX4 net5 A2 VSS VPW NHVT11LL_CKT W=0.225u L=40.00n
XX1 net5 A1 VSS VPW NHVT11LL_CKT W=0.225u L=40.00n
XX2 Z B VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX0 Z net5 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX5 net24 A2 VDD VNW PHVT11LL_CKT W=0.48u L=40.00n
XX6 net5 A1 net24 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX3 net36 B VDD VNW PHVT11LL_CKT W=0.85u L=40.00n
XX9 Z net5 net36 VNW PHVT11LL_CKT W=0.85u L=40.00n
.ENDS OA1B2V3_12TH40
.SUBCKT OA1B2V4_12TH40 A1 A2 B Z VDD VSS
XX4 net5 A2 VSS VPW NHVT11LL_CKT W=0.285u L=40.00n
XX1 net5 A1 VSS VPW NHVT11LL_CKT W=0.285u L=40.00n
XX2 Z B VSS VPW NHVT11LL_CKT W=0.57u L=40.00n
XX0 Z net5 VSS VPW NHVT11LL_CKT W=0.57u L=40.00n
XX5 net24 A2 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX6 net5 A1 net24 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX3 net36 B VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX9 Z net5 net36 VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS OA1B2V4_12TH40
.SUBCKT OA1B2V6_12TH40 A1 A2 B Z VDD VSS
XX4 net5 A2 VSS VPW NHVT11LL_CKT W=0.46u L=40.00n
XX1 net5 A1 VSS VPW NHVT11LL_CKT W=0.46u L=40.00n
XX2 Z B VSS VPW NHVT11LL_CKT W=0.855u L=40.00n
XX0 Z net5 VSS VPW NHVT11LL_CKT W=0.855u L=40.00n
XX5 net24 A2 VDD VNW PHVT11LL_CKT W=0.98u L=40.00n
XX6 net5 A1 net24 VNW PHVT11LL_CKT W=0.98u L=40.00n
XX3 net36 B VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX9 Z net5 net36 VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS OA1B2V6_12TH40
.SUBCKT OA1B2V8_12TH40 A1 A2 B Z VDD VSS
XX4 net5 A2 VSS VPW NHVT11LL_CKT W=0.645u L=40.00n
XX1 net5 A1 VSS VPW NHVT11LL_CKT W=0.645u L=40.00n
XX2 Z B VSS VPW NHVT11LL_CKT W=1.14u L=40.00n
XX0 Z net5 VSS VPW NHVT11LL_CKT W=1.14u L=40.00n
XX5 net24 A2 VDD VNW PHVT11LL_CKT W=1.38u L=40.00n
XX6 net5 A1 net24 VNW PHVT11LL_CKT W=1.38u L=40.00n
XX3 net36 B VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX9 Z net5 net36 VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS OA1B2V8_12TH40
.SUBCKT OA211V0_12TH40 A1 A2 B C Z VDD VSS
XX8 Z net18 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX0 net38 A2 VSS VPW NHVT11LL_CKT W=0.505u L=40.00n
XX2 net38 A1 VSS VPW NHVT11LL_CKT W=0.505u L=40.00n
XX5 net34 B net38 VPW NHVT11LL_CKT W=0.505u L=40.00n
XX6 net18 C net34 VPW NHVT11LL_CKT W=0.505u L=40.00n
XX1 net18 B VDD VNW PHVT11LL_CKT W=0.235u L=40.00n
XX7 Z net18 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX9 net18 A1 net21 VNW PHVT11LL_CKT W=0.44u L=40.00n
XX3 net21 A2 VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX4 net18 C VDD VNW PHVT11LL_CKT W=0.235u L=40.00n
.ENDS OA211V0_12TH40
.SUBCKT OA211V12_12TH40 A1 A2 B C Z VDD VSS
XX8 Z net18 VSS VPW NHVT11LL_CKT W=3.21u L=40.00n
XX0 net38 A2 VSS VPW NHVT11LL_CKT W=4.68u L=40.00n
XX2 net38 A1 VSS VPW NHVT11LL_CKT W=4.68u L=40.00n
XX5 net34 B net38 VPW NHVT11LL_CKT W=4.68u L=40.00n
XX6 net18 C net34 VPW NHVT11LL_CKT W=4.68u L=40.00n
XX1 net18 B VDD VNW PHVT11LL_CKT W=2.2u L=40.00n
XX7 Z net18 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX9 net18 A1 net21 VNW PHVT11LL_CKT W=4.12u L=40.00n
XX3 net21 A2 VDD VNW PHVT11LL_CKT W=4.12u L=40.00n
XX4 net18 C VDD VNW PHVT11LL_CKT W=2.2u L=40.00n
.ENDS OA211V12_12TH40
.SUBCKT OA211V1_12TH40 A1 A2 B C Z VDD VSS
XX8 Z net18 VSS VPW NHVT11LL_CKT W=0.375u L=40.00n
XX0 net38 A2 VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX2 net38 A1 VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX5 net34 B net38 VPW NHVT11LL_CKT W=0.61u L=40.00n
XX6 net18 C net34 VPW NHVT11LL_CKT W=0.61u L=40.00n
XX1 net18 B VDD VNW PHVT11LL_CKT W=0.285u L=40.00n
XX7 Z net18 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX9 net18 A1 net21 VNW PHVT11LL_CKT W=0.535u L=40.00n
XX3 net21 A2 VDD VNW PHVT11LL_CKT W=0.535u L=40.00n
XX4 net18 C VDD VNW PHVT11LL_CKT W=0.285u L=40.00n
.ENDS OA211V1_12TH40
.SUBCKT OA211V2_12TH40 A1 A2 B C Z VDD VSS
XX8 Z net18 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX0 net38 A2 VSS VPW NHVT11LL_CKT W=880.00n L=40.00n
XX2 net38 A1 VSS VPW NHVT11LL_CKT W=880.00n L=40.00n
XX5 net34 B net38 VPW NHVT11LL_CKT W=880.00n L=40.00n
XX6 net18 C net34 VPW NHVT11LL_CKT W=880.00n L=40.00n
XX1 net18 B VDD VNW PHVT11LL_CKT W=410.00n L=40.00n
XX7 Z net18 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX9 net18 A1 net21 VNW PHVT11LL_CKT W=770.00n L=40.00n
XX3 net21 A2 VDD VNW PHVT11LL_CKT W=770.00n L=40.00n
XX4 net18 C VDD VNW PHVT11LL_CKT W=410.00n L=40.00n
.ENDS OA211V2_12TH40
.SUBCKT OA211V3_12TH40 A1 A2 B C Z VDD VSS
XX8 Z net18 VSS VPW NHVT11LL_CKT W=0.75u L=40.00n
XX0 net38 A2 VSS VPW NHVT11LL_CKT W=1.14u L=40.00n
XX2 net38 A1 VSS VPW NHVT11LL_CKT W=1.14u L=40.00n
XX5 net34 B net38 VPW NHVT11LL_CKT W=1.14u L=40.00n
XX6 net18 C net34 VPW NHVT11LL_CKT W=1.14u L=40.00n
XX1 net18 B VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX7 Z net18 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX9 net18 A1 net21 VNW PHVT11LL_CKT W=1u L=40.00n
XX3 net21 A2 VDD VNW PHVT11LL_CKT W=1u L=40.00n
XX4 net18 C VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
.ENDS OA211V3_12TH40
.SUBCKT OA211V4_12TH40 A1 A2 B C Z VDD VSS
XX8 Z net18 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX0 net38 A2 VSS VPW NHVT11LL_CKT W=1.635u L=40.00n
XX2 net38 A1 VSS VPW NHVT11LL_CKT W=1.635u L=40.00n
XX5 net34 B net38 VPW NHVT11LL_CKT W=1.635u L=40.00n
XX6 net18 C net34 VPW NHVT11LL_CKT W=1.635u L=40.00n
XX1 net18 B VDD VNW PHVT11LL_CKT W=0.765u L=40.00n
XX7 Z net18 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX9 net18 A1 net21 VNW PHVT11LL_CKT W=1.44u L=40.00n
XX3 net21 A2 VDD VNW PHVT11LL_CKT W=1.44u L=40.00n
XX4 net18 C VDD VNW PHVT11LL_CKT W=0.765u L=40.00n
.ENDS OA211V4_12TH40
.SUBCKT OA211V6_12TH40 A1 A2 B C Z VDD VSS
XX8 Z net18 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX0 net38 A2 VSS VPW NHVT11LL_CKT W=2.32u L=40.00n
XX2 net38 A1 VSS VPW NHVT11LL_CKT W=2.32u L=40.00n
XX5 net34 B net38 VPW NHVT11LL_CKT W=2.32u L=40.00n
XX6 net18 C net34 VPW NHVT11LL_CKT W=2.32u L=40.00n
XX1 net18 B VDD VNW PHVT11LL_CKT W=1.1u L=40.00n
XX7 Z net18 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX9 net18 A1 net21 VNW PHVT11LL_CKT W=2.04u L=40.00n
XX3 net21 A2 VDD VNW PHVT11LL_CKT W=2.04u L=40.00n
XX4 net18 C VDD VNW PHVT11LL_CKT W=1.1u L=40.00n
.ENDS OA211V6_12TH40
.SUBCKT OA211V8_12TH40 A1 A2 B C Z VDD VSS
XX8 Z net18 VSS VPW NHVT11LL_CKT W=2.14u L=40.00n
XX0 net38 A2 VSS VPW NHVT11LL_CKT W=3.05u L=40.00n
XX2 net38 A1 VSS VPW NHVT11LL_CKT W=3.05u L=40.00n
XX5 net34 B net38 VPW NHVT11LL_CKT W=3.05u L=40.00n
XX6 net18 C net34 VPW NHVT11LL_CKT W=3.05u L=40.00n
XX1 net18 B VDD VNW PHVT11LL_CKT W=1.425u L=40.00n
XX7 Z net18 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX9 net18 A1 net21 VNW PHVT11LL_CKT W=2.675u L=40.00n
XX3 net21 A2 VDD VNW PHVT11LL_CKT W=2.675u L=40.00n
XX4 net18 C VDD VNW PHVT11LL_CKT W=1.425u L=40.00n
.ENDS OA211V8_12TH40
.SUBCKT OA21BV0_12TH40 A1 A2 B Z VDD VSS
XX6 net076 A2 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX11 Z B VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX10 Z net076 VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX5 net076 A1 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX4 net12 A2 VDD VNW PHVT11LL_CKT W=0.255u L=40.00n
XX1 net076 A1 net12 VNW PHVT11LL_CKT W=0.255u L=40.00n
XX8 net019 net076 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX9 Z B net019 VNW PHVT11LL_CKT W=0.305u L=40.00n
.ENDS OA21BV0_12TH40
.SUBCKT OA21BV12_12TH40 A1 A2 B Z VDD VSS
XX6 net076 A2 VSS VPW NHVT11LL_CKT W=0.855u L=40.00n
XX11 Z B VSS VPW NHVT11LL_CKT W=1.71u L=40.00n
XX10 Z net076 VSS VPW NHVT11LL_CKT W=1.71u L=40.00n
XX5 net076 A1 VSS VPW NHVT11LL_CKT W=0.855u L=40.00n
XX4 net12 A2 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX1 net076 A1 net12 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX8 net019 net076 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX9 Z B net019 VNW PHVT11LL_CKT W=3.66u L=40.00n
.ENDS OA21BV12_12TH40
.SUBCKT OA21BV16_12TH40 A1 A2 B Z VDD VSS
XX6 net076 A2 VSS VPW NHVT11LL_CKT W=1.35u L=40.00n
XX11 Z B VSS VPW NHVT11LL_CKT W=2.28u L=40.00n
XX10 Z net076 VSS VPW NHVT11LL_CKT W=2.28u L=40.00n
XX5 net076 A1 VSS VPW NHVT11LL_CKT W=1.35u L=40.00n
XX4 net12 A2 VDD VNW PHVT11LL_CKT W=2.9u L=40.00n
XX1 net076 A1 net12 VNW PHVT11LL_CKT W=2.9u L=40.00n
XX8 net019 net076 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX9 Z B net019 VNW PHVT11LL_CKT W=4.88u L=40.00n
.ENDS OA21BV16_12TH40
.SUBCKT OA21BV1_12TH40 A1 A2 B Z VDD VSS
XX6 net076 A2 VSS VPW NHVT11LL_CKT W=0.135u L=40.00n
XX11 Z B VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX10 Z net076 VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX5 net076 A1 VSS VPW NHVT11LL_CKT W=0.135u L=40.00n
XX4 net12 A2 VDD VNW PHVT11LL_CKT W=0.29u L=40.00n
XX1 net076 A1 net12 VNW PHVT11LL_CKT W=0.29u L=40.00n
XX8 net019 net076 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX9 Z B net019 VNW PHVT11LL_CKT W=0.43u L=40.00n
.ENDS OA21BV1_12TH40
.SUBCKT OA21BV2_12TH40 A1 A2 B Z VDD VSS
XX6 net076 A2 VSS VPW NHVT11LL_CKT W=170.00n L=40.00n
XX11 Z B VSS VPW NHVT11LL_CKT W=285.00n L=40.00n
XX10 Z net076 VSS VPW NHVT11LL_CKT W=285.00n L=40.00n
XX5 net076 A1 VSS VPW NHVT11LL_CKT W=170.00n L=40.00n
XX4 net12 A2 VDD VNW PHVT11LL_CKT W=365.00n L=40.00n
XX1 net076 A1 net12 VNW PHVT11LL_CKT W=365.00n L=40.00n
XX8 net019 net076 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX9 Z B net019 VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS OA21BV2_12TH40
.SUBCKT OA21BV3_12TH40 A1 A2 B Z VDD VSS
XX6 net076 A2 VSS VPW NHVT11LL_CKT W=0.225u L=40.00n
XX11 Z B VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX10 Z net076 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX5 net076 A1 VSS VPW NHVT11LL_CKT W=0.225u L=40.00n
XX4 net12 A2 VDD VNW PHVT11LL_CKT W=0.48u L=40.00n
XX1 net076 A1 net12 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX8 net019 net076 VDD VNW PHVT11LL_CKT W=0.85u L=40.00n
XX9 Z B net019 VNW PHVT11LL_CKT W=0.85u L=40.00n
.ENDS OA21BV3_12TH40
.SUBCKT OA21BV4_12TH40 A1 A2 B Z VDD VSS
XX6 net076 A2 VSS VPW NHVT11LL_CKT W=0.285u L=40.00n
XX11 Z B VSS VPW NHVT11LL_CKT W=0.57u L=40.00n
XX10 Z net076 VSS VPW NHVT11LL_CKT W=0.57u L=40.00n
XX5 net076 A1 VSS VPW NHVT11LL_CKT W=0.285u L=40.00n
XX4 net12 A2 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX1 net076 A1 net12 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX8 net019 net076 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX9 Z B net019 VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS OA21BV4_12TH40
.SUBCKT OA21BV6_12TH40 A1 A2 B Z VDD VSS
XX6 net076 A2 VSS VPW NHVT11LL_CKT W=0.46u L=40.00n
XX11 Z B VSS VPW NHVT11LL_CKT W=0.855u L=40.00n
XX10 Z net076 VSS VPW NHVT11LL_CKT W=0.855u L=40.00n
XX5 net076 A1 VSS VPW NHVT11LL_CKT W=0.46u L=40.00n
XX4 net12 A2 VDD VNW PHVT11LL_CKT W=0.98u L=40.00n
XX1 net076 A1 net12 VNW PHVT11LL_CKT W=0.98u L=40.00n
XX8 net019 net076 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX9 Z B net019 VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS OA21BV6_12TH40
.SUBCKT OA21BV8_12TH40 A1 A2 B Z VDD VSS
XX6 net076 A2 VSS VPW NHVT11LL_CKT W=0.645u L=40.00n
XX11 Z B VSS VPW NHVT11LL_CKT W=1.14u L=40.00n
XX10 Z net076 VSS VPW NHVT11LL_CKT W=1.14u L=40.00n
XX5 net076 A1 VSS VPW NHVT11LL_CKT W=0.645u L=40.00n
XX4 net12 A2 VDD VNW PHVT11LL_CKT W=1.38u L=40.00n
XX1 net076 A1 net12 VNW PHVT11LL_CKT W=1.38u L=40.00n
XX8 net019 net076 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX9 Z B net019 VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS OA21BV8_12TH40
.SUBCKT OA21V0_12TH40 A1 A2 B Z VDD VSS
XX5 net9 A1 VSS VPW NHVT11LL_CKT W=0.295u L=40.00n
XX6 net9 A2 VSS VPW NHVT11LL_CKT W=0.295u L=40.00n
XX8 net21 B net9 VPW NHVT11LL_CKT W=0.295u L=40.00n
XX0 Z net21 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX1 net21 A1 net24 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX4 net24 A2 VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX7 net21 B VDD VNW PHVT11LL_CKT W=0.195u L=40.00n
XX3 Z net21 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
.ENDS OA21V0_12TH40
.SUBCKT OA21V12_12TH40 A1 A2 B Z VDD VSS
XX5 net9 A1 VSS VPW NHVT11LL_CKT W=2.525u L=40.00n
XX6 net9 A2 VSS VPW NHVT11LL_CKT W=2.525u L=40.00n
XX8 net21 B net9 VPW NHVT11LL_CKT W=2.525u L=40.00n
XX0 Z net21 VSS VPW NHVT11LL_CKT W=3.21u L=40.00n
XX1 net21 A1 net24 VNW PHVT11LL_CKT W=3.05u L=40.00n
XX4 net24 A2 VDD VNW PHVT11LL_CKT W=3.05u L=40.00n
XX7 net21 B VDD VNW PHVT11LL_CKT W=1.625u L=40.00n
XX3 Z net21 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
.ENDS OA21V12_12TH40
.SUBCKT OA21V16_12TH40 A1 A2 B Z VDD VSS
XX5 net9 A1 VSS VPW NHVT11LL_CKT W=3.325u L=40.00n
XX6 net9 A2 VSS VPW NHVT11LL_CKT W=3.325u L=40.00n
XX8 net21 B net9 VPW NHVT11LL_CKT W=3.325u L=40.00n
XX0 Z net21 VSS VPW NHVT11LL_CKT W=4.28u L=40.00n
XX1 net21 A1 net24 VNW PHVT11LL_CKT W=4.025u L=40.00n
XX4 net24 A2 VDD VNW PHVT11LL_CKT W=4.025u L=40.00n
XX7 net21 B VDD VNW PHVT11LL_CKT W=2.17u L=40.00n
XX3 Z net21 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
.ENDS OA21V16_12TH40
.SUBCKT OA21V1_12TH40 A1 A2 B Z VDD VSS
XX5 net9 A1 VSS VPW NHVT11LL_CKT W=0.365u L=40.00n
XX6 net9 A2 VSS VPW NHVT11LL_CKT W=0.365u L=40.00n
XX8 net21 B net9 VPW NHVT11LL_CKT W=0.365u L=40.00n
XX0 Z net21 VSS VPW NHVT11LL_CKT W=0.375u L=40.00n
XX1 net21 A1 net24 VNW PHVT11LL_CKT W=0.44u L=40.00n
XX4 net24 A2 VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX7 net21 B VDD VNW PHVT11LL_CKT W=0.235u L=40.00n
XX3 Z net21 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
.ENDS OA21V1_12TH40
.SUBCKT OA21V2_12TH40 A1 A2 B Z VDD VSS
XX5 net9 A1 VSS VPW NHVT11LL_CKT W=465.00n L=40.00n
XX6 net9 A2 VSS VPW NHVT11LL_CKT W=465.00n L=40.00n
XX8 net21 B net9 VPW NHVT11LL_CKT W=465.00n L=40.00n
XX0 Z net21 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX1 net21 A1 net24 VNW PHVT11LL_CKT W=565.00n L=40.00n
XX4 net24 A2 VDD VNW PHVT11LL_CKT W=565.00n L=40.00n
XX7 net21 B VDD VNW PHVT11LL_CKT W=305.00n L=40.00n
XX3 Z net21 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS OA21V2_12TH40
.SUBCKT OA21V3_12TH40 A1 A2 B Z VDD VSS
XX5 net9 A1 VSS VPW NHVT11LL_CKT W=670.00n L=40.00n
XX6 net9 A2 VSS VPW NHVT11LL_CKT W=670.00n L=40.00n
XX8 net21 B net9 VPW NHVT11LL_CKT W=670.00n L=40.00n
XX0 Z net21 VSS VPW NHVT11LL_CKT W=0.75u L=40.00n
XX1 net21 A1 net24 VNW PHVT11LL_CKT W=810.00n L=40.00n
XX4 net24 A2 VDD VNW PHVT11LL_CKT W=810.00n L=40.00n
XX7 net21 B VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX3 Z net21 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
.ENDS OA21V3_12TH40
.SUBCKT OA21V4_12TH40 A1 A2 B Z VDD VSS
XX5 net9 A1 VSS VPW NHVT11LL_CKT W=870.00n L=40.00n
XX6 net9 A2 VSS VPW NHVT11LL_CKT W=870.00n L=40.00n
XX8 net21 B net9 VPW NHVT11LL_CKT W=870.00n L=40.00n
XX0 Z net21 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX1 net21 A1 net24 VNW PHVT11LL_CKT W=1.05u L=40.00n
XX4 net24 A2 VDD VNW PHVT11LL_CKT W=1.05u L=40.00n
XX7 net21 B VDD VNW PHVT11LL_CKT W=560.00n L=40.00n
XX3 Z net21 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS OA21V4_12TH40
.SUBCKT OA21V6_12TH40 A1 A2 B Z VDD VSS
XX5 net9 A1 VSS VPW NHVT11LL_CKT W=1.305u L=40.00n
XX6 net9 A2 VSS VPW NHVT11LL_CKT W=1.305u L=40.00n
XX8 net21 B net9 VPW NHVT11LL_CKT W=1.305u L=40.00n
XX0 Z net21 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX1 net21 A1 net24 VNW PHVT11LL_CKT W=1.575u L=40.00n
XX4 net24 A2 VDD VNW PHVT11LL_CKT W=1.575u L=40.00n
XX7 net21 B VDD VNW PHVT11LL_CKT W=0.84u L=40.00n
XX3 Z net21 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS OA21V6_12TH40
.SUBCKT OA21V8_12TH40 A1 A2 B Z VDD VSS
XX5 net9 A1 VSS VPW NHVT11LL_CKT W=1.7u L=40.00n
XX6 net9 A2 VSS VPW NHVT11LL_CKT W=1.7u L=40.00n
XX8 net21 B net9 VPW NHVT11LL_CKT W=1.7u L=40.00n
XX0 Z net21 VSS VPW NHVT11LL_CKT W=2.14u L=40.00n
XX1 net21 A1 net24 VNW PHVT11LL_CKT W=2.04u L=40.00n
XX4 net24 A2 VDD VNW PHVT11LL_CKT W=2.04u L=40.00n
XX7 net21 B VDD VNW PHVT11LL_CKT W=1.1u L=40.00n
XX3 Z net21 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS OA21V8_12TH40
.SUBCKT OA221V1_12TH40 A1 A2 B1 B2 C Z VDD VSS
XX8 net10 B2 net18 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX6 net060 C net10 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX5 net10 B1 net18 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX2 net18 A1 VSS VPW NHVT11LL_CKT W=430.00n L=40.00n
XX0 net18 A2 VSS VPW NHVT11LL_CKT W=430.00n L=40.00n
XX10 Z net060 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX11 Z net060 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX7 net060 B1 net084 VNW PHVT11LL_CKT W=380.00n L=40.00n
XX4 net060 C VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX3 net33 A2 VDD VNW PHVT11LL_CKT W=380.00n L=40.00n
XX9 net060 A1 net33 VNW PHVT11LL_CKT W=380.00n L=40.00n
XX1 net084 B2 VDD VNW PHVT11LL_CKT W=380.00n L=40.00n
.ENDS OA221V1_12TH40
.SUBCKT OA221V2_12TH40 A1 A2 B1 B2 C Z VDD VSS
XX8 net10 B2 net18 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX6 net060 C net10 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX5 net10 B1 net18 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX2 net18 A1 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX0 net18 A2 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX10 Z net060 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX11 Z net060 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX7 net060 B1 net084 VNW PHVT11LL_CKT W=540.00n L=40.00n
XX4 net060 C VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
XX3 net33 A2 VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX9 net060 A1 net33 VNW PHVT11LL_CKT W=540.00n L=40.00n
XX1 net084 B2 VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
.ENDS OA221V2_12TH40
.SUBCKT OA221V4_12TH40 A1 A2 B1 B2 C Z VDD VSS
XX8 net10 B2 net18 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX6 net060 C net10 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX5 net10 B1 net18 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX2 net18 A1 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX0 net18 A2 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX10 Z net060 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX11 Z net060 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX7 net060 B1 net084 VNW PHVT11LL_CKT W=1.08u L=40.00n
XX4 net060 C VDD VNW PHVT11LL_CKT W=620.00n L=40.00n
XX3 net33 A2 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX9 net060 A1 net33 VNW PHVT11LL_CKT W=1.08u L=40.00n
XX1 net084 B2 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
.ENDS OA221V4_12TH40
.SUBCKT OA221V8_12TH40 A1 A2 B1 B2 C Z VDD VSS
XX8 net10 B2 net18 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX6 net060 C net10 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX5 net10 B1 net18 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX2 net18 A1 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX0 net18 A2 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX10 Z net060 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX11 Z net060 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX7 net060 B1 net084 VNW PHVT11LL_CKT W=2.16u L=40.00n
XX4 net060 C VDD VNW PHVT11LL_CKT W=1.24u L=40.00n
XX3 net33 A2 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
XX9 net060 A1 net33 VNW PHVT11LL_CKT W=2.16u L=40.00n
XX1 net084 B2 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
.ENDS OA221V8_12TH40
.SUBCKT OA222V1_12TH40 A1 A2 B1 B2 C1 C2 Z VDD VSS
XX10 net065 C2 net52 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX12 Z net065 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX0 net40 A2 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX2 net40 A1 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX5 net52 B1 net40 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX6 net065 C1 net52 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX8 net52 B2 net40 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX13 Z net065 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX11 net065 C1 net11 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX1 net31 B2 VDD VNW PHVT11LL_CKT W=0.38u L=40.00n
XX9 net065 A1 net23 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX3 net23 A2 VDD VNW PHVT11LL_CKT W=0.38u L=40.00n
XX4 net11 C2 VDD VNW PHVT11LL_CKT W=0.38u L=40.00n
XX7 net065 B1 net31 VNW PHVT11LL_CKT W=0.38u L=40.00n
.ENDS OA222V1_12TH40
.SUBCKT OA222V2_12TH40 A1 A2 B1 B2 C1 C2 Z VDD VSS
XX10 net065 C2 net52 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX12 Z net065 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX0 net40 A2 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX2 net40 A1 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX5 net52 B1 net40 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX6 net065 C1 net52 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX8 net52 B2 net40 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX13 Z net065 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX11 net065 C1 net11 VNW PHVT11LL_CKT W=540.00n L=40.00n
XX1 net31 B2 VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX9 net065 A1 net23 VNW PHVT11LL_CKT W=540.00n L=40.00n
XX3 net23 A2 VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX4 net11 C2 VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX7 net065 B1 net31 VNW PHVT11LL_CKT W=540.00n L=40.00n
.ENDS OA222V2_12TH40
.SUBCKT OA222V4_12TH40 A1 A2 B1 B2 C1 C2 Z VDD VSS
XX10 net065 C2 net52 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX12 Z net065 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX0 net40 A2 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX2 net40 A1 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX5 net52 B1 net40 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX6 net065 C1 net52 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX8 net52 B2 net40 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX13 Z net065 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX11 net065 C1 net11 VNW PHVT11LL_CKT W=1.08u L=40.00n
XX1 net31 B2 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX9 net065 A1 net23 VNW PHVT11LL_CKT W=1.08u L=40.00n
XX3 net23 A2 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX4 net11 C2 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX7 net065 B1 net31 VNW PHVT11LL_CKT W=1.08u L=40.00n
.ENDS OA222V4_12TH40
.SUBCKT OA222V8_12TH40 A1 A2 B1 B2 C1 C2 Z VDD VSS
XX10 net065 C2 net52 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX12 Z net065 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX0 net40 A2 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX2 net40 A1 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX5 net52 B1 net40 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX6 net065 C1 net52 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX8 net52 B2 net40 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX13 Z net065 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX11 net065 C1 net11 VNW PHVT11LL_CKT W=2.16u L=40.00n
XX1 net31 B2 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
XX9 net065 A1 net23 VNW PHVT11LL_CKT W=2.16u L=40.00n
XX3 net23 A2 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
XX4 net11 C2 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
XX7 net065 B1 net31 VNW PHVT11LL_CKT W=2.16u L=40.00n
.ENDS OA222V8_12TH40
.SUBCKT OA22V0_12TH40 A1 A2 B1 B2 Z VDD VSS
XX9 net30 B2 net38 VPW NHVT11LL_CKT W=0.31u L=40.00n
XX0 Z net30 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX8 net30 B1 net38 VPW NHVT11LL_CKT W=0.31u L=40.00n
XX6 net38 A2 VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX5 net38 A1 VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX2 net13 B2 VDD VNW PHVT11LL_CKT W=0.37u L=40.00n
XX3 Z net30 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX7 net30 B1 net13 VNW PHVT11LL_CKT W=0.37u L=40.00n
XX4 net25 A2 VDD VNW PHVT11LL_CKT W=0.37u L=40.00n
XX1 net30 A1 net25 VNW PHVT11LL_CKT W=0.37u L=40.00n
.ENDS OA22V0_12TH40
.SUBCKT OA22V12_12TH40 A1 A2 B1 B2 Z VDD VSS
XX9 net30 B2 net38 VPW NHVT11LL_CKT W=2.79u L=40.00n
XX0 Z net30 VSS VPW NHVT11LL_CKT W=3.21u L=40.00n
XX8 net30 B1 net38 VPW NHVT11LL_CKT W=2.79u L=40.00n
XX6 net38 A2 VSS VPW NHVT11LL_CKT W=2.79u L=40.00n
XX5 net38 A1 VSS VPW NHVT11LL_CKT W=2.79u L=40.00n
XX2 net13 B2 VDD VNW PHVT11LL_CKT W=3.36u L=40.00n
XX3 Z net30 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX7 net30 B1 net13 VNW PHVT11LL_CKT W=3.36u L=40.00n
XX4 net25 A2 VDD VNW PHVT11LL_CKT W=3.36u L=40.00n
XX1 net30 A1 net25 VNW PHVT11LL_CKT W=3.36u L=40.00n
.ENDS OA22V12_12TH40
.SUBCKT OA22V16_12TH40 A1 A2 B1 B2 Z VDD VSS
XX9 net30 B2 net38 VPW NHVT11LL_CKT W=3.72u L=40.00n
XX0 Z net30 VSS VPW NHVT11LL_CKT W=4.28u L=40.00n
XX8 net30 B1 net38 VPW NHVT11LL_CKT W=3.72u L=40.00n
XX6 net38 A2 VSS VPW NHVT11LL_CKT W=3.72u L=40.00n
XX5 net38 A1 VSS VPW NHVT11LL_CKT W=3.72u L=40.00n
XX2 net13 B2 VDD VNW PHVT11LL_CKT W=4.52u L=40.00n
XX3 Z net30 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX7 net30 B1 net13 VNW PHVT11LL_CKT W=4.52u L=40.00n
XX4 net25 A2 VDD VNW PHVT11LL_CKT W=4.52u L=40.00n
XX1 net30 A1 net25 VNW PHVT11LL_CKT W=4.52u L=40.00n
.ENDS OA22V16_12TH40
.SUBCKT OA22V1_12TH40 A1 A2 B1 B2 Z VDD VSS
XX9 net30 B2 net38 VPW NHVT11LL_CKT W=0.375u L=40.00n
XX0 Z net30 VSS VPW NHVT11LL_CKT W=0.375u L=40.00n
XX8 net30 B1 net38 VPW NHVT11LL_CKT W=0.375u L=40.00n
XX6 net38 A2 VSS VPW NHVT11LL_CKT W=0.375u L=40.00n
XX5 net38 A1 VSS VPW NHVT11LL_CKT W=0.375u L=40.00n
XX2 net13 B2 VDD VNW PHVT11LL_CKT W=0.455u L=40.00n
XX3 Z net30 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX7 net30 B1 net13 VNW PHVT11LL_CKT W=0.455u L=40.00n
XX4 net25 A2 VDD VNW PHVT11LL_CKT W=0.455u L=40.00n
XX1 net30 A1 net25 VNW PHVT11LL_CKT W=0.455u L=40.00n
.ENDS OA22V1_12TH40
.SUBCKT OA22V2_12TH40 A1 A2 B1 B2 Z VDD VSS
XX9 net30 B2 net38 VPW NHVT11LL_CKT W=480.00n L=40.00n
XX0 Z net30 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX8 net30 B1 net38 VPW NHVT11LL_CKT W=480.00n L=40.00n
XX6 net38 A2 VSS VPW NHVT11LL_CKT W=480.00n L=40.00n
XX5 net38 A1 VSS VPW NHVT11LL_CKT W=480.00n L=40.00n
XX2 net13 B2 VDD VNW PHVT11LL_CKT W=580.00n L=40.00n
XX3 Z net30 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX7 net30 B1 net13 VNW PHVT11LL_CKT W=580.00n L=40.00n
XX4 net25 A2 VDD VNW PHVT11LL_CKT W=580.00n L=40.00n
XX1 net30 A1 net25 VNW PHVT11LL_CKT W=580.00n L=40.00n
.ENDS OA22V2_12TH40
.SUBCKT OA22V3_12TH40 A1 A2 B1 B2 Z VDD VSS
XX9 net30 B2 net38 VPW NHVT11LL_CKT W=0.75u L=40.00n
XX0 Z net30 VSS VPW NHVT11LL_CKT W=0.75u L=40.00n
XX8 net30 B1 net38 VPW NHVT11LL_CKT W=0.75u L=40.00n
XX6 net38 A2 VSS VPW NHVT11LL_CKT W=0.75u L=40.00n
XX5 net38 A1 VSS VPW NHVT11LL_CKT W=0.75u L=40.00n
XX2 net13 B2 VDD VNW PHVT11LL_CKT W=0.9u L=40.00n
XX3 Z net30 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX7 net30 B1 net13 VNW PHVT11LL_CKT W=0.9u L=40.00n
XX4 net25 A2 VDD VNW PHVT11LL_CKT W=0.9u L=40.00n
XX1 net30 A1 net25 VNW PHVT11LL_CKT W=0.9u L=40.00n
.ENDS OA22V3_12TH40
.SUBCKT OA22V4_12TH40 A1 A2 B1 B2 Z VDD VSS
XX9 net30 B2 net38 VPW NHVT11LL_CKT W=0.95u L=40.00n
XX0 Z net30 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX8 net30 B1 net38 VPW NHVT11LL_CKT W=0.95u L=40.00n
XX6 net38 A2 VSS VPW NHVT11LL_CKT W=0.95u L=40.00n
XX5 net38 A1 VSS VPW NHVT11LL_CKT W=0.95u L=40.00n
XX2 net13 B2 VDD VNW PHVT11LL_CKT W=1.15u L=40.00n
XX3 Z net30 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX7 net30 B1 net13 VNW PHVT11LL_CKT W=1.15u L=40.00n
XX4 net25 A2 VDD VNW PHVT11LL_CKT W=1.15u L=40.00n
XX1 net30 A1 net25 VNW PHVT11LL_CKT W=1.15u L=40.00n
.ENDS OA22V4_12TH40
.SUBCKT OA22V6_12TH40 A1 A2 B1 B2 Z VDD VSS
XX9 net30 B2 net38 VPW NHVT11LL_CKT W=1.47u L=40.00n
XX0 Z net30 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX8 net30 B1 net38 VPW NHVT11LL_CKT W=1.47u L=40.00n
XX6 net38 A2 VSS VPW NHVT11LL_CKT W=1.47u L=40.00n
XX5 net38 A1 VSS VPW NHVT11LL_CKT W=1.47u L=40.00n
XX2 net13 B2 VDD VNW PHVT11LL_CKT W=1.77u L=40.00n
XX3 Z net30 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX7 net30 B1 net13 VNW PHVT11LL_CKT W=1.77u L=40.00n
XX4 net25 A2 VDD VNW PHVT11LL_CKT W=1.77u L=40.00n
XX1 net30 A1 net25 VNW PHVT11LL_CKT W=1.77u L=40.00n
.ENDS OA22V6_12TH40
.SUBCKT OA22V8_12TH40 A1 A2 B1 B2 Z VDD VSS
XX9 net30 B2 net38 VPW NHVT11LL_CKT W=1.88u L=40.00n
XX0 Z net30 VSS VPW NHVT11LL_CKT W=2.14u L=40.00n
XX8 net30 B1 net38 VPW NHVT11LL_CKT W=1.88u L=40.00n
XX6 net38 A2 VSS VPW NHVT11LL_CKT W=1.88u L=40.00n
XX5 net38 A1 VSS VPW NHVT11LL_CKT W=1.88u L=40.00n
XX2 net13 B2 VDD VNW PHVT11LL_CKT W=2.28u L=40.00n
XX3 Z net30 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX7 net30 B1 net13 VNW PHVT11LL_CKT W=2.28u L=40.00n
XX4 net25 A2 VDD VNW PHVT11LL_CKT W=2.28u L=40.00n
XX1 net30 A1 net25 VNW PHVT11LL_CKT W=2.28u L=40.00n
.ENDS OA22V8_12TH40
.SUBCKT OA31V1_12TH40 A1 A2 A3 B Z VDD VSS
XX2 net6 A3 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX5 net6 A1 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX6 net6 A2 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX8 net047 B net6 VPW NHVT11LL_CKT W=250.00n L=40.00n
XX4 Z net047 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX9 Z net047 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX3 net29 A3 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX0 net33 A2 net29 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX7 net047 A1 net33 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX1 net047 B VDD VNW PHVT11LL_CKT W=180.00n L=40.00n
.ENDS OA31V1_12TH40
.SUBCKT OA31V2_12TH40 A1 A2 A3 B Z VDD VSS
XX2 net6 A3 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX5 net6 A1 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX6 net6 A2 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX8 net047 B net6 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX4 Z net047 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX9 Z net047 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX3 net29 A3 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX0 net33 A2 net29 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX7 net047 A1 net33 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 net047 B VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
.ENDS OA31V2_12TH40
.SUBCKT OA31V4_12TH40 A1 A2 A3 B Z VDD VSS
XX2 net6 A3 VSS VPW NHVT11LL_CKT W=700.00n L=40.00n
XX5 net6 A1 VSS VPW NHVT11LL_CKT W=700.00n L=40.00n
XX6 net6 A2 VSS VPW NHVT11LL_CKT W=700.00n L=40.00n
XX8 net047 B net6 VPW NHVT11LL_CKT W=700.00n L=40.00n
XX4 Z net047 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX9 Z net047 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX3 net29 A3 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 net33 A2 net29 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX7 net047 A1 net33 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 net047 B VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
.ENDS OA31V4_12TH40
.SUBCKT OA31V8_12TH40 A1 A2 A3 B Z VDD VSS
XX2 net6 A3 VSS VPW NHVT11LL_CKT W=1.4u L=40.00n
XX5 net6 A1 VSS VPW NHVT11LL_CKT W=1.4u L=40.00n
XX6 net6 A2 VSS VPW NHVT11LL_CKT W=1.4u L=40.00n
XX8 net047 B net6 VPW NHVT11LL_CKT W=1.4u L=40.00n
XX4 Z net047 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX9 Z net047 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX3 net29 A3 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX0 net33 A2 net29 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX7 net047 A1 net33 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 net047 B VDD VNW PHVT11LL_CKT W=1.00u L=40.00n
.ENDS OA31V8_12TH40
.SUBCKT OA32V1_12TH40 A1 A2 A3 B1 B2 Z VDD VSS
XX10 Z net022 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX9 net022 B2 net6 VPW NHVT11LL_CKT W=250.00n L=40.00n
XX2 net6 A3 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX5 net6 A1 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX6 net6 A2 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX8 net022 B1 net6 VPW NHVT11LL_CKT W=250.00n L=40.00n
XX11 Z net022 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX4 net055 B2 VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
XX3 net29 A3 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX0 net33 A2 net29 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX7 net022 A1 net33 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX1 net022 B1 net055 VNW PHVT11LL_CKT W=310.00n L=40.00n
.ENDS OA32V1_12TH40
.SUBCKT OA32V2_12TH40 A1 A2 A3 B1 B2 Z VDD VSS
XX10 Z net022 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX9 net022 B2 net6 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX2 net6 A3 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX5 net6 A1 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX6 net6 A2 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX8 net022 B1 net6 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX11 Z net022 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX4 net055 B2 VDD VNW PHVT11LL_CKT W=460.00n L=40.00n
XX3 net29 A3 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX0 net33 A2 net29 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX7 net022 A1 net33 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 net022 B1 net055 VNW PHVT11LL_CKT W=460.00n L=40.00n
.ENDS OA32V2_12TH40
.SUBCKT OA32V4_12TH40 A1 A2 A3 B1 B2 Z VDD VSS
XX10 Z net022 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX9 net022 B2 net6 VPW NHVT11LL_CKT W=700.00n L=40.00n
XX2 net6 A3 VSS VPW NHVT11LL_CKT W=700.00n L=40.00n
XX5 net6 A1 VSS VPW NHVT11LL_CKT W=700.00n L=40.00n
XX6 net6 A2 VSS VPW NHVT11LL_CKT W=700.00n L=40.00n
XX8 net022 B1 net6 VPW NHVT11LL_CKT W=700.00n L=40.00n
XX11 Z net022 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX4 net055 B2 VDD VNW PHVT11LL_CKT W=920.00n L=40.00n
XX3 net29 A3 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 net33 A2 net29 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX7 net022 A1 net33 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 net022 B1 net055 VNW PHVT11LL_CKT W=920.00n L=40.00n
.ENDS OA32V4_12TH40
.SUBCKT OA32V8_12TH40 A1 A2 A3 B1 B2 Z VDD VSS
XX10 Z net022 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX9 net022 B2 net6 VPW NHVT11LL_CKT W=1.4u L=40.00n
XX2 net6 A3 VSS VPW NHVT11LL_CKT W=1.4u L=40.00n
XX5 net6 A1 VSS VPW NHVT11LL_CKT W=1.4u L=40.00n
XX6 net6 A2 VSS VPW NHVT11LL_CKT W=1.4u L=40.00n
XX8 net022 B1 net6 VPW NHVT11LL_CKT W=1.4u L=40.00n
XX11 Z net022 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX4 net055 B2 VDD VNW PHVT11LL_CKT W=1.84u L=40.00n
XX3 net29 A3 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX0 net33 A2 net29 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX7 net022 A1 net33 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 net022 B1 net055 VNW PHVT11LL_CKT W=1.84u L=40.00n
.ENDS OA32V8_12TH40
.SUBCKT OA33V1_12TH40 A1 A2 A3 B1 B2 B3 Z VDD VSS
XX12 Z net025 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX11 net025 B3 net6 VPW NHVT11LL_CKT W=250.00n L=40.00n
XX9 net025 B2 net6 VPW NHVT11LL_CKT W=250.00n L=40.00n
XX2 net6 A3 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX5 net6 A1 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX6 net6 A2 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX8 net025 B1 net6 VPW NHVT11LL_CKT W=250.00n L=40.00n
XX13 Z net025 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX10 net050 B3 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX4 net055 B2 net050 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX3 net29 A3 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX0 net33 A2 net29 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX7 net025 A1 net33 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX1 net025 B1 net055 VNW PHVT11LL_CKT W=430.00n L=40.00n
.ENDS OA33V1_12TH40
.SUBCKT OA33V2_12TH40 A1 A2 A3 B1 B2 B3 Z VDD VSS
XX12 Z net025 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX11 net025 B3 net6 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX9 net025 B2 net6 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX2 net6 A3 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX5 net6 A1 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX6 net6 A2 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX8 net025 B1 net6 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX13 Z net025 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX10 net050 B3 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX4 net055 B2 net050 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX3 net29 A3 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX0 net33 A2 net29 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX7 net025 A1 net33 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 net025 B1 net055 VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS OA33V2_12TH40
.SUBCKT OA33V4_12TH40 A1 A2 A3 B1 B2 B3 Z VDD VSS
XX12 Z net025 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX11 net025 B3 net6 VPW NHVT11LL_CKT W=700.00n L=40.00n
XX9 net025 B2 net6 VPW NHVT11LL_CKT W=700.00n L=40.00n
XX2 net6 A3 VSS VPW NHVT11LL_CKT W=700.00n L=40.00n
XX5 net6 A1 VSS VPW NHVT11LL_CKT W=700.00n L=40.00n
XX6 net6 A2 VSS VPW NHVT11LL_CKT W=700.00n L=40.00n
XX8 net025 B1 net6 VPW NHVT11LL_CKT W=700.00n L=40.00n
XX13 Z net025 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX10 net050 B3 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX4 net055 B2 net050 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX3 net29 A3 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 net33 A2 net29 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX7 net025 A1 net33 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 net025 B1 net055 VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS OA33V4_12TH40
.SUBCKT OA33V8_12TH40 A1 A2 A3 B1 B2 B3 Z VDD VSS
XX12 Z net025 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX11 net025 B3 net6 VPW NHVT11LL_CKT W=1.4u L=40.00n
XX9 net025 B2 net6 VPW NHVT11LL_CKT W=1.4u L=40.00n
XX2 net6 A3 VSS VPW NHVT11LL_CKT W=1.4u L=40.00n
XX5 net6 A1 VSS VPW NHVT11LL_CKT W=1.4u L=40.00n
XX6 net6 A2 VSS VPW NHVT11LL_CKT W=1.4u L=40.00n
XX8 net025 B1 net6 VPW NHVT11LL_CKT W=1.4u L=40.00n
XX13 Z net025 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX10 net050 B3 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX4 net055 B2 net050 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX3 net29 A3 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX0 net33 A2 net29 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX7 net025 A1 net33 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 net025 B1 net055 VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS OA33V8_12TH40
.SUBCKT OAI211V0_12TH40 A1 A2 B C ZN VDD VSS
XX9 ZN C net34 VPW NHVT11LL_CKT W=0.295u L=40.00n
XX8 net34 B net38 VPW NHVT11LL_CKT W=0.295u L=40.00n
XX6 net38 A2 VSS VPW NHVT11LL_CKT W=0.295u L=40.00n
XX5 net38 A1 VSS VPW NHVT11LL_CKT W=0.295u L=40.00n
XX2 ZN C VDD VNW PHVT11LL_CKT W=0.13u L=40.00n
XX7 ZN B VDD VNW PHVT11LL_CKT W=0.13u L=40.00n
XX4 net25 A2 VDD VNW PHVT11LL_CKT W=0.255u L=40.00n
XX1 ZN A1 net25 VNW PHVT11LL_CKT W=0.255u L=40.00n
.ENDS OAI211V0_12TH40
.SUBCKT OAI211V1_12TH40 A1 A2 B C ZN VDD VSS
XX9 ZN C net34 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX8 net34 B net38 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX6 net38 A2 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX5 net38 A1 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX2 ZN C VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX7 ZN B VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX4 net25 A2 VDD VNW PHVT11LL_CKT W=0.375u L=40.00n
XX1 ZN A1 net25 VNW PHVT11LL_CKT W=0.375u L=40.00n
.ENDS OAI211V1_12TH40
.SUBCKT OAI211V2_12TH40 A1 A2 B C ZN VDD VSS
XX9 ZN C net34 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX8 net34 B net38 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX6 net38 A2 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX5 net38 A1 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX2 ZN C VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX7 ZN B VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX4 net25 A2 VDD VNW PHVT11LL_CKT W=535.00n L=40.00n
XX1 ZN A1 net25 VNW PHVT11LL_CKT W=535.00n L=40.00n
.ENDS OAI211V2_12TH40
.SUBCKT OAI211V3_12TH40 A1 A2 B C ZN VDD VSS
XX9 ZN C net34 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX8 net34 B net38 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX6 net38 A2 VSS VPW NHVT11LL_CKT W=0.86u L=40.00n
XX5 net38 A1 VSS VPW NHVT11LL_CKT W=0.86u L=40.00n
XX2 ZN C VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX7 ZN B VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX4 net25 A2 VDD VNW PHVT11LL_CKT W=0.75u L=40.00n
XX1 ZN A1 net25 VNW PHVT11LL_CKT W=0.75u L=40.00n
.ENDS OAI211V3_12TH40
.SUBCKT OAI211V4_12TH40 A1 A2 B C ZN VDD VSS
XX9 ZN C net34 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX8 net34 B net38 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX6 net38 A2 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX5 net38 A1 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX2 ZN C VDD VNW PHVT11LL_CKT W=0.57u L=40.00n
XX7 ZN B VDD VNW PHVT11LL_CKT W=0.57u L=40.00n
XX4 net25 A2 VDD VNW PHVT11LL_CKT W=1.07u L=40.00n
XX1 ZN A1 net25 VNW PHVT11LL_CKT W=1.07u L=40.00n
.ENDS OAI211V4_12TH40
.SUBCKT OAI211V6_12TH40 A1 A2 B C ZN VDD VSS
XX9 ZN C net34 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX8 net34 B net38 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX6 net38 A2 VSS VPW NHVT11LL_CKT W=1.83u L=40.00n
XX5 net38 A1 VSS VPW NHVT11LL_CKT W=1.83u L=40.00n
XX2 ZN C VDD VNW PHVT11LL_CKT W=0.855u L=40.00n
XX7 ZN B VDD VNW PHVT11LL_CKT W=0.855u L=40.00n
XX4 net25 A2 VDD VNW PHVT11LL_CKT W=1.605u L=40.00n
XX1 ZN A1 net25 VNW PHVT11LL_CKT W=1.605u L=40.00n
.ENDS OAI211V6_12TH40
.SUBCKT OAI211V8_12TH40 A1 A2 B C ZN VDD VSS
XX9 ZN C net34 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX8 net34 B net38 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX6 net38 A2 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX5 net38 A1 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX2 ZN C VDD VNW PHVT11LL_CKT W=1.14u L=40.00n
XX7 ZN B VDD VNW PHVT11LL_CKT W=1.14u L=40.00n
XX4 net25 A2 VDD VNW PHVT11LL_CKT W=2.14u L=40.00n
XX1 ZN A1 net25 VNW PHVT11LL_CKT W=2.14u L=40.00n
.ENDS OAI211V8_12TH40
.SUBCKT OAI21BV0_12TH40 A B1 B2 ZN VDD VSS
XX0 net21 A VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX8 ZN net21 net29 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX6 net29 B2 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX5 net29 B1 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX3 net21 A VDD VNW PHVT11LL_CKT W=0.135u L=40.00n
XX7 ZN net21 VDD VNW PHVT11LL_CKT W=0.165u L=40.00n
XX4 net20 B2 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX1 ZN B1 net20 VNW PHVT11LL_CKT W=0.305u L=40.00n
.ENDS OAI21BV0_12TH40
.SUBCKT OAI21BV12_12TH40 A B1 B2 ZN VDD VSS
XX0 net21 A VSS VPW NHVT11LL_CKT W=0.67u L=40.00n
XX8 ZN net21 net29 VPW NHVT11LL_CKT W=3.03u L=40.00n
XX6 net29 B2 VSS VPW NHVT11LL_CKT W=3.03u L=40.00n
XX5 net29 B1 VSS VPW NHVT11LL_CKT W=3.03u L=40.00n
XX3 net21 A VDD VNW PHVT11LL_CKT W=0.77u L=40.00n
XX7 ZN net21 VDD VNW PHVT11LL_CKT W=1.95u L=40.00n
XX4 net20 B2 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX1 ZN B1 net20 VNW PHVT11LL_CKT W=3.66u L=40.00n
.ENDS OAI21BV12_12TH40
.SUBCKT OAI21BV16_12TH40 A B1 B2 ZN VDD VSS
XX0 net21 A VSS VPW NHVT11LL_CKT W=0.89u L=40.00n
XX8 ZN net21 net29 VPW NHVT11LL_CKT W=4.04u L=40.00n
XX6 net29 B2 VSS VPW NHVT11LL_CKT W=4.04u L=40.00n
XX5 net29 B1 VSS VPW NHVT11LL_CKT W=4.04u L=40.00n
XX3 net21 A VDD VNW PHVT11LL_CKT W=1.01u L=40.00n
XX7 ZN net21 VDD VNW PHVT11LL_CKT W=2.6u L=40.00n
XX4 net20 B2 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX1 ZN B1 net20 VNW PHVT11LL_CKT W=4.88u L=40.00n
.ENDS OAI21BV16_12TH40
.SUBCKT OAI21BV1_12TH40 A B1 B2 ZN VDD VSS
XX0 net21 A VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX8 ZN net21 net29 VPW NHVT11LL_CKT W=0.355u L=40.00n
XX6 net29 B2 VSS VPW NHVT11LL_CKT W=0.355u L=40.00n
XX5 net29 B1 VSS VPW NHVT11LL_CKT W=0.355u L=40.00n
XX3 net21 A VDD VNW PHVT11LL_CKT W=0.135u L=40.00n
XX7 ZN net21 VDD VNW PHVT11LL_CKT W=0.23u L=40.00n
XX4 net20 B2 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX1 ZN B1 net20 VNW PHVT11LL_CKT W=0.43u L=40.00n
.ENDS OAI21BV1_12TH40
.SUBCKT OAI21BV2_12TH40 A B1 B2 ZN VDD VSS
XX0 net21 A VSS VPW NHVT11LL_CKT W=135.00n L=40.00n
XX8 ZN net21 net29 VPW NHVT11LL_CKT W=505.00n L=40.00n
XX6 net29 B2 VSS VPW NHVT11LL_CKT W=505.00n L=40.00n
XX5 net29 B1 VSS VPW NHVT11LL_CKT W=505.00n L=40.00n
XX3 net21 A VDD VNW PHVT11LL_CKT W=155.00n L=40.00n
XX7 ZN net21 VDD VNW PHVT11LL_CKT W=325.00n L=40.00n
XX4 net20 B2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 ZN B1 net20 VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS OAI21BV2_12TH40
.SUBCKT OAI21BV3_12TH40 A B1 B2 ZN VDD VSS
XX0 net21 A VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX8 ZN net21 net29 VPW NHVT11LL_CKT W=0.71u L=40.00n
XX6 net29 B2 VSS VPW NHVT11LL_CKT W=0.71u L=40.00n
XX5 net29 B1 VSS VPW NHVT11LL_CKT W=0.71u L=40.00n
XX3 net21 A VDD VNW PHVT11LL_CKT W=0.205u L=40.00n
XX7 ZN net21 VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
XX4 net20 B2 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX1 ZN B1 net20 VNW PHVT11LL_CKT W=0.86u L=40.00n
.ENDS OAI21BV3_12TH40
.SUBCKT OAI21BV4_12TH40 A B1 B2 ZN VDD VSS
XX0 net21 A VSS VPW NHVT11LL_CKT W=0.24u L=40.00n
XX8 ZN net21 net29 VPW NHVT11LL_CKT W=1.01u L=40.00n
XX6 net29 B2 VSS VPW NHVT11LL_CKT W=1.01u L=40.00n
XX5 net29 B1 VSS VPW NHVT11LL_CKT W=1.01u L=40.00n
XX3 net21 A VDD VNW PHVT11LL_CKT W=0.27u L=40.00n
XX7 ZN net21 VDD VNW PHVT11LL_CKT W=0.65u L=40.00n
XX4 net20 B2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 ZN B1 net20 VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS OAI21BV4_12TH40
.SUBCKT OAI21BV6_12TH40 A B1 B2 ZN VDD VSS
XX0 net21 A VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX8 ZN net21 net29 VPW NHVT11LL_CKT W=1.515u L=40.00n
XX6 net29 B2 VSS VPW NHVT11LL_CKT W=1.515u L=40.00n
XX5 net29 B1 VSS VPW NHVT11LL_CKT W=1.515u L=40.00n
XX3 net21 A VDD VNW PHVT11LL_CKT W=0.39u L=40.00n
XX7 ZN net21 VDD VNW PHVT11LL_CKT W=0.975u L=40.00n
XX4 net20 B2 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX1 ZN B1 net20 VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS OAI21BV6_12TH40
.SUBCKT OAI21BV8_12TH40 A B1 B2 ZN VDD VSS
XX0 net21 A VSS VPW NHVT11LL_CKT W=0.45u L=40.00n
XX8 ZN net21 net29 VPW NHVT11LL_CKT W=2.02u L=40.00n
XX6 net29 B2 VSS VPW NHVT11LL_CKT W=2.02u L=40.00n
XX5 net29 B1 VSS VPW NHVT11LL_CKT W=2.02u L=40.00n
XX3 net21 A VDD VNW PHVT11LL_CKT W=0.51u L=40.00n
XX7 ZN net21 VDD VNW PHVT11LL_CKT W=1.3u L=40.00n
XX4 net20 B2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 ZN B1 net20 VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS OAI21BV8_12TH40
.SUBCKT OAI21V0_12TH40 A1 A2 B ZN VDD VSS
XX8 ZN B net29 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX6 net29 A2 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX5 net29 A1 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX7 ZN B VDD VNW PHVT11LL_CKT W=0.165u L=40.00n
XX4 net20 A2 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX1 ZN A1 net20 VNW PHVT11LL_CKT W=0.305u L=40.00n
.ENDS OAI21V0_12TH40
.SUBCKT OAI21V12_12TH40 A1 A2 B ZN VDD VSS
XX8 ZN B net29 VPW NHVT11LL_CKT W=3.03u L=40.00n
XX6 net29 A2 VSS VPW NHVT11LL_CKT W=3.03u L=40.00n
XX5 net29 A1 VSS VPW NHVT11LL_CKT W=3.03u L=40.00n
XX7 ZN B VDD VNW PHVT11LL_CKT W=1.95u L=40.00n
XX4 net20 A2 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX1 ZN A1 net20 VNW PHVT11LL_CKT W=3.66u L=40.00n
.ENDS OAI21V12_12TH40
.SUBCKT OAI21V16_12TH40 A1 A2 B ZN VDD VSS
XX8 ZN B net29 VPW NHVT11LL_CKT W=4.04u L=40.00n
XX6 net29 A2 VSS VPW NHVT11LL_CKT W=4.04u L=40.00n
XX5 net29 A1 VSS VPW NHVT11LL_CKT W=4.04u L=40.00n
XX7 ZN B VDD VNW PHVT11LL_CKT W=2.6u L=40.00n
XX4 net20 A2 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX1 ZN A1 net20 VNW PHVT11LL_CKT W=4.88u L=40.00n
.ENDS OAI21V16_12TH40
.SUBCKT OAI21V1_12TH40 A1 A2 B ZN VDD VSS
XX8 ZN B net29 VPW NHVT11LL_CKT W=0.355u L=40.00n
XX6 net29 A2 VSS VPW NHVT11LL_CKT W=0.355u L=40.00n
XX5 net29 A1 VSS VPW NHVT11LL_CKT W=0.355u L=40.00n
XX7 ZN B VDD VNW PHVT11LL_CKT W=0.23u L=40.00n
XX4 net20 A2 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX1 ZN A1 net20 VNW PHVT11LL_CKT W=0.43u L=40.00n
.ENDS OAI21V1_12TH40
.SUBCKT OAI21V2_12TH40 A1 A2 B ZN VDD VSS
XX8 ZN B net29 VPW NHVT11LL_CKT W=505.00n L=40.00n
XX6 net29 A2 VSS VPW NHVT11LL_CKT W=505.00n L=40.00n
XX5 net29 A1 VSS VPW NHVT11LL_CKT W=505.00n L=40.00n
XX7 ZN B VDD VNW PHVT11LL_CKT W=325.00n L=40.00n
XX4 net20 A2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 ZN A1 net20 VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS OAI21V2_12TH40
.SUBCKT OAI21V3_12TH40 A1 A2 B ZN VDD VSS
XX8 ZN B net29 VPW NHVT11LL_CKT W=0.71u L=40.00n
XX6 net29 A2 VSS VPW NHVT11LL_CKT W=0.71u L=40.00n
XX5 net29 A1 VSS VPW NHVT11LL_CKT W=0.71u L=40.00n
XX7 ZN B VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
XX4 net20 A2 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX1 ZN A1 net20 VNW PHVT11LL_CKT W=0.86u L=40.00n
.ENDS OAI21V3_12TH40
.SUBCKT OAI21V4_12TH40 A1 A2 B ZN VDD VSS
XX8 ZN B net29 VPW NHVT11LL_CKT W=1.01u L=40.00n
XX6 net29 A2 VSS VPW NHVT11LL_CKT W=1.01u L=40.00n
XX5 net29 A1 VSS VPW NHVT11LL_CKT W=1.01u L=40.00n
XX7 ZN B VDD VNW PHVT11LL_CKT W=0.65u L=40.00n
XX4 net20 A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 ZN A1 net20 VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS OAI21V4_12TH40
.SUBCKT OAI21V6_12TH40 A1 A2 B ZN VDD VSS
XX8 ZN B net29 VPW NHVT11LL_CKT W=1.515u L=40.00n
XX6 net29 A2 VSS VPW NHVT11LL_CKT W=1.515u L=40.00n
XX5 net29 A1 VSS VPW NHVT11LL_CKT W=1.515u L=40.00n
XX7 ZN B VDD VNW PHVT11LL_CKT W=0.975u L=40.00n
XX4 net20 A2 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX1 ZN A1 net20 VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS OAI21V6_12TH40
.SUBCKT OAI21V8_12TH40 A1 A2 B ZN VDD VSS
XX8 ZN B net29 VPW NHVT11LL_CKT W=2.02u L=40.00n
XX6 net29 A2 VSS VPW NHVT11LL_CKT W=2.02u L=40.00n
XX5 net29 A1 VSS VPW NHVT11LL_CKT W=2.02u L=40.00n
XX7 ZN B VDD VNW PHVT11LL_CKT W=1.3u L=40.00n
XX4 net20 A2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 ZN A1 net20 VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS OAI21V8_12TH40
.SUBCKT OAI221V0_12TH40 A1 A2 B1 B2 C ZN VDD VSS
XX8 net10 B2 net18 VPW NHVT11LL_CKT W=0.305u L=40.00n
XX6 ZN C net10 VPW NHVT11LL_CKT W=0.305u L=40.00n
XX5 net10 B1 net18 VPW NHVT11LL_CKT W=0.305u L=40.00n
XX2 net18 A1 VSS VPW NHVT11LL_CKT W=0.305u L=40.00n
XX0 net18 A2 VSS VPW NHVT11LL_CKT W=0.305u L=40.00n
XX7 ZN B1 net084 VNW PHVT11LL_CKT W=0.265u L=40.00n
XX4 ZN C VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX3 net33 A2 VDD VNW PHVT11LL_CKT W=0.265u L=40.00n
XX9 ZN A1 net33 VNW PHVT11LL_CKT W=0.265u L=40.00n
XX1 net084 B2 VDD VNW PHVT11LL_CKT W=0.265u L=40.00n
.ENDS OAI221V0_12TH40
.SUBCKT OAI221V1_12TH40 A1 A2 B1 B2 C ZN VDD VSS
XX8 net10 B2 net18 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX6 ZN C net10 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX5 net10 B1 net18 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX2 net18 A1 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX0 net18 A2 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX7 ZN B1 net084 VNW PHVT11LL_CKT W=0.375u L=40.00n
XX4 ZN C VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX3 net33 A2 VDD VNW PHVT11LL_CKT W=0.375u L=40.00n
XX9 ZN A1 net33 VNW PHVT11LL_CKT W=0.375u L=40.00n
XX1 net084 B2 VDD VNW PHVT11LL_CKT W=0.375u L=40.00n
.ENDS OAI221V1_12TH40
.SUBCKT OAI221V2_12TH40 A1 A2 B1 B2 C ZN VDD VSS
XX8 net10 B2 net18 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX6 ZN C net10 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX5 net10 B1 net18 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX2 net18 A1 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX0 net18 A2 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX7 ZN B1 net084 VNW PHVT11LL_CKT W=535.00n L=40.00n
XX4 ZN C VDD VNW PHVT11LL_CKT W=285.00n L=40.00n
XX3 net33 A2 VDD VNW PHVT11LL_CKT W=535.00n L=40.00n
XX9 ZN A1 net33 VNW PHVT11LL_CKT W=535.00n L=40.00n
XX1 net084 B2 VDD VNW PHVT11LL_CKT W=535.00n L=40.00n
.ENDS OAI221V2_12TH40
.SUBCKT OAI221V3_12TH40 A1 A2 B1 B2 C ZN VDD VSS
XX8 net10 B2 net18 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX6 ZN C net10 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX5 net10 B1 net18 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX2 net18 A1 VSS VPW NHVT11LL_CKT W=0.86u L=40.00n
XX0 net18 A2 VSS VPW NHVT11LL_CKT W=0.86u L=40.00n
XX7 ZN B1 net084 VNW PHVT11LL_CKT W=0.75u L=40.00n
XX4 ZN C VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX3 net33 A2 VDD VNW PHVT11LL_CKT W=0.75u L=40.00n
XX9 ZN A1 net33 VNW PHVT11LL_CKT W=0.75u L=40.00n
XX1 net084 B2 VDD VNW PHVT11LL_CKT W=0.75u L=40.00n
.ENDS OAI221V3_12TH40
.SUBCKT OAI221V4_12TH40 A1 A2 B1 B2 C ZN VDD VSS
XX8 net10 B2 net18 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX6 ZN C net10 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX5 net10 B1 net18 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX2 net18 A1 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX0 net18 A2 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX7 ZN B1 net084 VNW PHVT11LL_CKT W=1.07u L=40.00n
XX4 ZN C VDD VNW PHVT11LL_CKT W=0.57u L=40.00n
XX3 net33 A2 VDD VNW PHVT11LL_CKT W=1.07u L=40.00n
XX9 ZN A1 net33 VNW PHVT11LL_CKT W=1.07u L=40.00n
XX1 net084 B2 VDD VNW PHVT11LL_CKT W=1.07u L=40.00n
.ENDS OAI221V4_12TH40
.SUBCKT OAI221V6_12TH40 A1 A2 B1 B2 C ZN VDD VSS
XX8 net10 B2 net18 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX6 ZN C net10 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX5 net10 B1 net18 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX2 net18 A1 VSS VPW NHVT11LL_CKT W=1.83u L=40.00n
XX0 net18 A2 VSS VPW NHVT11LL_CKT W=1.83u L=40.00n
XX7 ZN B1 net084 VNW PHVT11LL_CKT W=1.605u L=40.00n
XX4 ZN C VDD VNW PHVT11LL_CKT W=0.855u L=40.00n
XX3 net33 A2 VDD VNW PHVT11LL_CKT W=1.605u L=40.00n
XX9 ZN A1 net33 VNW PHVT11LL_CKT W=1.605u L=40.00n
XX1 net084 B2 VDD VNW PHVT11LL_CKT W=1.605u L=40.00n
.ENDS OAI221V6_12TH40
.SUBCKT OAI221V8_12TH40 A1 A2 B1 B2 C ZN VDD VSS
XX8 net10 B2 net18 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX6 ZN C net10 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX5 net10 B1 net18 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX2 net18 A1 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX0 net18 A2 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX7 ZN B1 net084 VNW PHVT11LL_CKT W=2.14u L=40.00n
XX4 ZN C VDD VNW PHVT11LL_CKT W=1.14u L=40.00n
XX3 net33 A2 VDD VNW PHVT11LL_CKT W=2.14u L=40.00n
XX9 ZN A1 net33 VNW PHVT11LL_CKT W=2.14u L=40.00n
XX1 net084 B2 VDD VNW PHVT11LL_CKT W=2.14u L=40.00n
.ENDS OAI221V8_12TH40
.SUBCKT OAI222V0_12TH40 A1 A2 B1 B2 C1 C2 ZN VDD VSS
XX10 ZN C2 net52 VPW NHVT11LL_CKT W=0.305u L=40.00n
XX0 net40 A2 VSS VPW NHVT11LL_CKT W=0.305u L=40.00n
XX2 net40 A1 VSS VPW NHVT11LL_CKT W=0.305u L=40.00n
XX5 net52 B1 net40 VPW NHVT11LL_CKT W=0.305u L=40.00n
XX6 ZN C1 net52 VPW NHVT11LL_CKT W=0.305u L=40.00n
XX8 net52 B2 net40 VPW NHVT11LL_CKT W=0.305u L=40.00n
XX11 ZN C1 net11 VNW PHVT11LL_CKT W=0.265u L=40.00n
XX1 net31 B2 VDD VNW PHVT11LL_CKT W=0.265u L=40.00n
XX9 ZN A1 net23 VNW PHVT11LL_CKT W=0.265u L=40.00n
XX3 net23 A2 VDD VNW PHVT11LL_CKT W=0.265u L=40.00n
XX4 net11 C2 VDD VNW PHVT11LL_CKT W=0.265u L=40.00n
XX7 ZN B1 net31 VNW PHVT11LL_CKT W=0.265u L=40.00n
.ENDS OAI222V0_12TH40
.SUBCKT OAI222V1_12TH40 A1 A2 B1 B2 C1 C2 ZN VDD VSS
XX10 ZN C2 net52 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX0 net40 A2 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX2 net40 A1 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX5 net52 B1 net40 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX6 ZN C1 net52 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX8 net52 B2 net40 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX11 ZN C1 net11 VNW PHVT11LL_CKT W=0.375u L=40.00n
XX1 net31 B2 VDD VNW PHVT11LL_CKT W=0.375u L=40.00n
XX9 ZN A1 net23 VNW PHVT11LL_CKT W=0.375u L=40.00n
XX3 net23 A2 VDD VNW PHVT11LL_CKT W=0.375u L=40.00n
XX4 net11 C2 VDD VNW PHVT11LL_CKT W=0.375u L=40.00n
XX7 ZN B1 net31 VNW PHVT11LL_CKT W=0.375u L=40.00n
.ENDS OAI222V1_12TH40
.SUBCKT OAI222V2_12TH40 A1 A2 B1 B2 C1 C2 ZN VDD VSS
XX10 ZN C2 net52 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX0 net40 A2 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX2 net40 A1 VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX5 net52 B1 net40 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX6 ZN C1 net52 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX8 net52 B2 net40 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX11 ZN C1 net11 VNW PHVT11LL_CKT W=535.00n L=40.00n
XX1 net31 B2 VDD VNW PHVT11LL_CKT W=535.00n L=40.00n
XX9 ZN A1 net23 VNW PHVT11LL_CKT W=535.00n L=40.00n
XX3 net23 A2 VDD VNW PHVT11LL_CKT W=535.00n L=40.00n
XX4 net11 C2 VDD VNW PHVT11LL_CKT W=535.00n L=40.00n
XX7 ZN B1 net31 VNW PHVT11LL_CKT W=535.00n L=40.00n
.ENDS OAI222V2_12TH40
.SUBCKT OAI222V3_12TH40 A1 A2 B1 B2 C1 C2 ZN VDD VSS
XX10 ZN C2 net52 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX0 net40 A2 VSS VPW NHVT11LL_CKT W=0.86u L=40.00n
XX2 net40 A1 VSS VPW NHVT11LL_CKT W=0.86u L=40.00n
XX5 net52 B1 net40 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX6 ZN C1 net52 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX8 net52 B2 net40 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX11 ZN C1 net11 VNW PHVT11LL_CKT W=0.75u L=40.00n
XX1 net31 B2 VDD VNW PHVT11LL_CKT W=0.75u L=40.00n
XX9 ZN A1 net23 VNW PHVT11LL_CKT W=0.75u L=40.00n
XX3 net23 A2 VDD VNW PHVT11LL_CKT W=0.75u L=40.00n
XX4 net11 C2 VDD VNW PHVT11LL_CKT W=0.75u L=40.00n
XX7 ZN B1 net31 VNW PHVT11LL_CKT W=0.75u L=40.00n
.ENDS OAI222V3_12TH40
.SUBCKT OAI222V4_12TH40 A1 A2 B1 B2 C1 C2 ZN VDD VSS
XX10 ZN C2 net52 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX0 net40 A2 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX2 net40 A1 VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX5 net52 B1 net40 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX6 ZN C1 net52 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX8 net52 B2 net40 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX11 ZN C1 net11 VNW PHVT11LL_CKT W=1.07u L=40.00n
XX1 net31 B2 VDD VNW PHVT11LL_CKT W=1.07u L=40.00n
XX9 ZN A1 net23 VNW PHVT11LL_CKT W=1.07u L=40.00n
XX3 net23 A2 VDD VNW PHVT11LL_CKT W=1.07u L=40.00n
XX4 net11 C2 VDD VNW PHVT11LL_CKT W=1.07u L=40.00n
XX7 ZN B1 net31 VNW PHVT11LL_CKT W=1.07u L=40.00n
.ENDS OAI222V4_12TH40
.SUBCKT OAI222V6_12TH40 A1 A2 B1 B2 C1 C2 ZN VDD VSS
XX10 ZN C2 net52 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX0 net40 A2 VSS VPW NHVT11LL_CKT W=1.83u L=40.00n
XX2 net40 A1 VSS VPW NHVT11LL_CKT W=1.83u L=40.00n
XX5 net52 B1 net40 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX6 ZN C1 net52 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX8 net52 B2 net40 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX11 ZN C1 net11 VNW PHVT11LL_CKT W=1.605u L=40.00n
XX1 net31 B2 VDD VNW PHVT11LL_CKT W=1.605u L=40.00n
XX9 ZN A1 net23 VNW PHVT11LL_CKT W=1.605u L=40.00n
XX3 net23 A2 VDD VNW PHVT11LL_CKT W=1.605u L=40.00n
XX4 net11 C2 VDD VNW PHVT11LL_CKT W=1.605u L=40.00n
XX7 ZN B1 net31 VNW PHVT11LL_CKT W=1.605u L=40.00n
.ENDS OAI222V6_12TH40
.SUBCKT OAI222V8_12TH40 A1 A2 B1 B2 C1 C2 ZN VDD VSS
XX10 ZN C2 net52 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX0 net40 A2 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX2 net40 A1 VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX5 net52 B1 net40 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX6 ZN C1 net52 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX8 net52 B2 net40 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX11 ZN C1 net11 VNW PHVT11LL_CKT W=2.14u L=40.00n
XX1 net31 B2 VDD VNW PHVT11LL_CKT W=2.14u L=40.00n
XX9 ZN A1 net23 VNW PHVT11LL_CKT W=2.14u L=40.00n
XX3 net23 A2 VDD VNW PHVT11LL_CKT W=2.14u L=40.00n
XX4 net11 C2 VDD VNW PHVT11LL_CKT W=2.14u L=40.00n
XX7 ZN B1 net31 VNW PHVT11LL_CKT W=2.14u L=40.00n
.ENDS OAI222V8_12TH40
.SUBCKT OAI22BBV0_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX11 net26 A2 VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX8 ZN net10 net38 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX6 net38 B2 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX5 net38 B1 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX9 net10 A1 net26 VPW NHVT11LL_CKT W=0.185u L=40.00n
XX10 net10 A1 VDD VNW PHVT11LL_CKT W=0.125u L=40.00n
XX2 net10 A2 VDD VNW PHVT11LL_CKT W=0.125u L=40.00n
XX7 ZN net10 VDD VNW PHVT11LL_CKT W=0.165u L=40.00n
XX4 net25 B2 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX1 ZN B1 net25 VNW PHVT11LL_CKT W=0.305u L=40.00n
.ENDS OAI22BBV0_12TH40
.SUBCKT OAI22BBV12_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX11 net26 A2 VSS VPW NHVT11LL_CKT W=1.59u L=40.00n
XX8 ZN net10 net38 VPW NHVT11LL_CKT W=3.03u L=40.00n
XX6 net38 B2 VSS VPW NHVT11LL_CKT W=3.03u L=40.00n
XX5 net38 B1 VSS VPW NHVT11LL_CKT W=3.03u L=40.00n
XX9 net10 A1 net26 VPW NHVT11LL_CKT W=1.59u L=40.00n
XX10 net10 A1 VDD VNW PHVT11LL_CKT W=1.02u L=40.00n
XX2 net10 A2 VDD VNW PHVT11LL_CKT W=1.02u L=40.00n
XX7 ZN net10 VDD VNW PHVT11LL_CKT W=1.95u L=40.00n
XX4 net25 B2 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX1 ZN B1 net25 VNW PHVT11LL_CKT W=3.66u L=40.00n
.ENDS OAI22BBV12_12TH40
.SUBCKT OAI22BBV16_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX11 net26 A2 VSS VPW NHVT11LL_CKT W=2.06u L=40.00n
XX8 ZN net10 net38 VPW NHVT11LL_CKT W=4.04u L=40.00n
XX6 net38 B2 VSS VPW NHVT11LL_CKT W=4.04u L=40.00n
XX5 net38 B1 VSS VPW NHVT11LL_CKT W=4.04u L=40.00n
XX9 net10 A1 net26 VPW NHVT11LL_CKT W=2.06u L=40.00n
XX10 net10 A1 VDD VNW PHVT11LL_CKT W=1.34u L=40.00n
XX2 net10 A2 VDD VNW PHVT11LL_CKT W=1.34u L=40.00n
XX7 ZN net10 VDD VNW PHVT11LL_CKT W=2.6u L=40.00n
XX4 net25 B2 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX1 ZN B1 net25 VNW PHVT11LL_CKT W=4.88u L=40.00n
.ENDS OAI22BBV16_12TH40
.SUBCKT OAI22BBV1_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX11 net26 A2 VSS VPW NHVT11LL_CKT W=0.235u L=40.00n
XX8 ZN net10 net38 VPW NHVT11LL_CKT W=0.355u L=40.00n
XX6 net38 B2 VSS VPW NHVT11LL_CKT W=0.355u L=40.00n
XX5 net38 B1 VSS VPW NHVT11LL_CKT W=0.355u L=40.00n
XX9 net10 A1 net26 VPW NHVT11LL_CKT W=0.235u L=40.00n
XX10 net10 A1 VDD VNW PHVT11LL_CKT W=0.155u L=40.00n
XX2 net10 A2 VDD VNW PHVT11LL_CKT W=0.155u L=40.00n
XX7 ZN net10 VDD VNW PHVT11LL_CKT W=0.23u L=40.00n
XX4 net25 B2 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX1 ZN B1 net25 VNW PHVT11LL_CKT W=0.43u L=40.00n
.ENDS OAI22BBV1_12TH40
.SUBCKT OAI22BBV2_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX11 net26 A2 VSS VPW NHVT11LL_CKT W=295.00n L=40.00n
XX8 ZN net10 net38 VPW NHVT11LL_CKT W=505.00n L=40.00n
XX6 net38 B2 VSS VPW NHVT11LL_CKT W=505.00n L=40.00n
XX5 net38 B1 VSS VPW NHVT11LL_CKT W=505.00n L=40.00n
XX9 net10 A1 net26 VPW NHVT11LL_CKT W=295.00n L=40.00n
XX10 net10 A1 VDD VNW PHVT11LL_CKT W=190.00n L=40.00n
XX2 net10 A2 VDD VNW PHVT11LL_CKT W=190.00n L=40.00n
XX7 ZN net10 VDD VNW PHVT11LL_CKT W=325.00n L=40.00n
XX4 net25 B2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 ZN B1 net25 VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS OAI22BBV2_12TH40
.SUBCKT OAI22BBV3_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX11 net26 A2 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX8 ZN net10 net38 VPW NHVT11LL_CKT W=0.71u L=40.00n
XX6 net38 B2 VSS VPW NHVT11LL_CKT W=0.71u L=40.00n
XX5 net38 B1 VSS VPW NHVT11LL_CKT W=0.71u L=40.00n
XX9 net10 A1 net26 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX10 net10 A1 VDD VNW PHVT11LL_CKT W=0.255u L=40.00n
XX2 net10 A2 VDD VNW PHVT11LL_CKT W=0.255u L=40.00n
XX7 ZN net10 VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
XX4 net25 B2 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX1 ZN B1 net25 VNW PHVT11LL_CKT W=0.86u L=40.00n
.ENDS OAI22BBV3_12TH40
.SUBCKT OAI22BBV4_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX11 net26 A2 VSS VPW NHVT11LL_CKT W=0.525u L=40.00n
XX8 ZN net10 net38 VPW NHVT11LL_CKT W=1.01u L=40.00n
XX6 net38 B2 VSS VPW NHVT11LL_CKT W=1.01u L=40.00n
XX5 net38 B1 VSS VPW NHVT11LL_CKT W=1.01u L=40.00n
XX9 net10 A1 net26 VPW NHVT11LL_CKT W=0.525u L=40.00n
XX10 net10 A1 VDD VNW PHVT11LL_CKT W=0.335u L=40.00n
XX2 net10 A2 VDD VNW PHVT11LL_CKT W=0.335u L=40.00n
XX7 ZN net10 VDD VNW PHVT11LL_CKT W=0.65u L=40.00n
XX4 net25 B2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 ZN B1 net25 VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS OAI22BBV4_12TH40
.SUBCKT OAI22BBV6_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX11 net26 A2 VSS VPW NHVT11LL_CKT W=0.77u L=40.00n
XX8 ZN net10 net38 VPW NHVT11LL_CKT W=1.515u L=40.00n
XX6 net38 B2 VSS VPW NHVT11LL_CKT W=1.515u L=40.00n
XX5 net38 B1 VSS VPW NHVT11LL_CKT W=1.515u L=40.00n
XX9 net10 A1 net26 VPW NHVT11LL_CKT W=0.77u L=40.00n
XX10 net10 A1 VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX2 net10 A2 VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX7 ZN net10 VDD VNW PHVT11LL_CKT W=0.975u L=40.00n
XX4 net25 B2 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX1 ZN B1 net25 VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS OAI22BBV6_12TH40
.SUBCKT OAI22BBV8_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX11 net26 A2 VSS VPW NHVT11LL_CKT W=1.04u L=40.00n
XX8 ZN net10 net38 VPW NHVT11LL_CKT W=2.02u L=40.00n
XX6 net38 B2 VSS VPW NHVT11LL_CKT W=2.02u L=40.00n
XX5 net38 B1 VSS VPW NHVT11LL_CKT W=2.02u L=40.00n
XX9 net10 A1 net26 VPW NHVT11LL_CKT W=1.04u L=40.00n
XX10 net10 A1 VDD VNW PHVT11LL_CKT W=0.67u L=40.00n
XX2 net10 A2 VDD VNW PHVT11LL_CKT W=0.67u L=40.00n
XX7 ZN net10 VDD VNW PHVT11LL_CKT W=1.3u L=40.00n
XX4 net25 B2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 ZN B1 net25 VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS OAI22BBV8_12TH40
.SUBCKT OAI22V0_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX2 ZN B2 net18 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX5 net18 A1 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX6 net18 A2 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX8 ZN B1 net18 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX0 net37 B2 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX1 ZN A1 net29 VNW PHVT11LL_CKT W=0.305u L=40.00n
XX4 net29 A2 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX7 ZN B1 net37 VNW PHVT11LL_CKT W=0.305u L=40.00n
.ENDS OAI22V0_12TH40
.SUBCKT OAI22V12_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX2 ZN B2 net18 VPW NHVT11LL_CKT W=3.03u L=40.00n
XX5 net18 A1 VSS VPW NHVT11LL_CKT W=3.03u L=40.00n
XX6 net18 A2 VSS VPW NHVT11LL_CKT W=3.03u L=40.00n
XX8 ZN B1 net18 VPW NHVT11LL_CKT W=3.03u L=40.00n
XX0 net37 B2 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX1 ZN A1 net29 VNW PHVT11LL_CKT W=3.66u L=40.00n
XX4 net29 A2 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX7 ZN B1 net37 VNW PHVT11LL_CKT W=3.66u L=40.00n
.ENDS OAI22V12_12TH40
.SUBCKT OAI22V16_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX2 ZN B2 net18 VPW NHVT11LL_CKT W=4.04u L=40.00n
XX5 net18 A1 VSS VPW NHVT11LL_CKT W=4.04u L=40.00n
XX6 net18 A2 VSS VPW NHVT11LL_CKT W=4.04u L=40.00n
XX8 ZN B1 net18 VPW NHVT11LL_CKT W=4.04u L=40.00n
XX0 net37 B2 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX1 ZN A1 net29 VNW PHVT11LL_CKT W=4.88u L=40.00n
XX4 net29 A2 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX7 ZN B1 net37 VNW PHVT11LL_CKT W=4.88u L=40.00n
.ENDS OAI22V16_12TH40
.SUBCKT OAI22V1_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX2 ZN B2 net18 VPW NHVT11LL_CKT W=0.355u L=40.00n
XX5 net18 A1 VSS VPW NHVT11LL_CKT W=0.355u L=40.00n
XX6 net18 A2 VSS VPW NHVT11LL_CKT W=0.355u L=40.00n
XX8 ZN B1 net18 VPW NHVT11LL_CKT W=0.355u L=40.00n
XX0 net37 B2 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX1 ZN A1 net29 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX4 net29 A2 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX7 ZN B1 net37 VNW PHVT11LL_CKT W=0.43u L=40.00n
.ENDS OAI22V1_12TH40
.SUBCKT OAI22V2_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX2 ZN B2 net18 VPW NHVT11LL_CKT W=505.00n L=40.00n
XX5 net18 A1 VSS VPW NHVT11LL_CKT W=505.00n L=40.00n
XX6 net18 A2 VSS VPW NHVT11LL_CKT W=505.00n L=40.00n
XX8 ZN B1 net18 VPW NHVT11LL_CKT W=505.00n L=40.00n
XX0 net37 B2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 ZN A1 net29 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX4 net29 A2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX7 ZN B1 net37 VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS OAI22V2_12TH40
.SUBCKT OAI22V3_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX2 ZN B2 net18 VPW NHVT11LL_CKT W=0.71u L=40.00n
XX5 net18 A1 VSS VPW NHVT11LL_CKT W=0.71u L=40.00n
XX6 net18 A2 VSS VPW NHVT11LL_CKT W=0.71u L=40.00n
XX8 ZN B1 net18 VPW NHVT11LL_CKT W=0.71u L=40.00n
XX0 net37 B2 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX1 ZN A1 net29 VNW PHVT11LL_CKT W=0.86u L=40.00n
XX4 net29 A2 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX7 ZN B1 net37 VNW PHVT11LL_CKT W=0.86u L=40.00n
.ENDS OAI22V3_12TH40
.SUBCKT OAI22V4_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX2 ZN B2 net18 VPW NHVT11LL_CKT W=1.01u L=40.00n
XX5 net18 A1 VSS VPW NHVT11LL_CKT W=1.01u L=40.00n
XX6 net18 A2 VSS VPW NHVT11LL_CKT W=1.01u L=40.00n
XX8 ZN B1 net18 VPW NHVT11LL_CKT W=1.01u L=40.00n
XX0 net37 B2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 ZN A1 net29 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX4 net29 A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX7 ZN B1 net37 VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS OAI22V4_12TH40
.SUBCKT OAI22V6_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX2 ZN B2 net18 VPW NHVT11LL_CKT W=1.515u L=40.00n
XX5 net18 A1 VSS VPW NHVT11LL_CKT W=1.515u L=40.00n
XX6 net18 A2 VSS VPW NHVT11LL_CKT W=1.515u L=40.00n
XX8 ZN B1 net18 VPW NHVT11LL_CKT W=1.515u L=40.00n
XX0 net37 B2 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX1 ZN A1 net29 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX4 net29 A2 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX7 ZN B1 net37 VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS OAI22V6_12TH40
.SUBCKT OAI22V8_12TH40 A1 A2 B1 B2 ZN VDD VSS
XX2 ZN B2 net18 VPW NHVT11LL_CKT W=2.02u L=40.00n
XX5 net18 A1 VSS VPW NHVT11LL_CKT W=2.02u L=40.00n
XX6 net18 A2 VSS VPW NHVT11LL_CKT W=2.02u L=40.00n
XX8 ZN B1 net18 VPW NHVT11LL_CKT W=2.02u L=40.00n
XX0 net37 B2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 ZN A1 net29 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX4 net29 A2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX7 ZN B1 net37 VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS OAI22V8_12TH40
.SUBCKT OAI2XB1V0_12TH40 A B1 B2 ZN VDD VSS
XX3 net21 B2 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX6 net29 net21 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX5 net29 B1 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX8 ZN A net29 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX2 net21 B2 VDD VNW PHVT11LL_CKT W=0.135u L=40.00n
XX7 ZN B1 net16 VNW PHVT11LL_CKT W=0.305u L=40.00n
XX1 ZN A VDD VNW PHVT11LL_CKT W=0.165u L=40.00n
XX0 net16 net21 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
.ENDS OAI2XB1V0_12TH40
.SUBCKT OAI2XB1V12_12TH40 A B1 B2 ZN VDD VSS
XX3 net21 B2 VSS VPW NHVT11LL_CKT W=0.87u L=40.00n
XX6 net29 net21 VSS VPW NHVT11LL_CKT W=3.03u L=40.00n
XX5 net29 B1 VSS VPW NHVT11LL_CKT W=3.03u L=40.00n
XX8 ZN A net29 VPW NHVT11LL_CKT W=3.03u L=40.00n
XX2 net21 B2 VDD VNW PHVT11LL_CKT W=1u L=40.00n
XX7 ZN B1 net16 VNW PHVT11LL_CKT W=3.66u L=40.00n
XX1 ZN A VDD VNW PHVT11LL_CKT W=1.95u L=40.00n
XX0 net16 net21 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
.ENDS OAI2XB1V12_12TH40
.SUBCKT OAI2XB1V16_12TH40 A B1 B2 ZN VDD VSS
XX3 net21 B2 VSS VPW NHVT11LL_CKT W=1.185u L=40.00n
XX6 net29 net21 VSS VPW NHVT11LL_CKT W=4.04u L=40.00n
XX5 net29 B1 VSS VPW NHVT11LL_CKT W=4.04u L=40.00n
XX8 ZN A net29 VPW NHVT11LL_CKT W=4.04u L=40.00n
XX2 net21 B2 VDD VNW PHVT11LL_CKT W=1.35u L=40.00n
XX7 ZN B1 net16 VNW PHVT11LL_CKT W=4.88u L=40.00n
XX1 ZN A VDD VNW PHVT11LL_CKT W=2.6u L=40.00n
XX0 net16 net21 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
.ENDS OAI2XB1V16_12TH40
.SUBCKT OAI2XB1V1_12TH40 A B1 B2 ZN VDD VSS
XX3 net21 B2 VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX6 net29 net21 VSS VPW NHVT11LL_CKT W=0.355u L=40.00n
XX5 net29 B1 VSS VPW NHVT11LL_CKT W=0.355u L=40.00n
XX8 ZN A net29 VPW NHVT11LL_CKT W=0.355u L=40.00n
XX2 net21 B2 VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX7 ZN B1 net16 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX1 ZN A VDD VNW PHVT11LL_CKT W=0.23u L=40.00n
XX0 net16 net21 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
.ENDS OAI2XB1V1_12TH40
.SUBCKT OAI2XB1V2_12TH40 A B1 B2 ZN VDD VSS
XX3 net21 B2 VSS VPW NHVT11LL_CKT W=170.00n L=40.00n
XX6 net29 net21 VSS VPW NHVT11LL_CKT W=505.00n L=40.00n
XX5 net29 B1 VSS VPW NHVT11LL_CKT W=505.00n L=40.00n
XX8 ZN A net29 VPW NHVT11LL_CKT W=505.00n L=40.00n
XX2 net21 B2 VDD VNW PHVT11LL_CKT W=195.00n L=40.00n
XX7 ZN B1 net16 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 ZN A VDD VNW PHVT11LL_CKT W=325.00n L=40.00n
XX0 net16 net21 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS OAI2XB1V2_12TH40
.SUBCKT OAI2XB1V3_12TH40 A B1 B2 ZN VDD VSS
XX3 net21 B2 VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX6 net29 net21 VSS VPW NHVT11LL_CKT W=0.71u L=40.00n
XX5 net29 B1 VSS VPW NHVT11LL_CKT W=0.71u L=40.00n
XX8 ZN A net29 VPW NHVT11LL_CKT W=0.71u L=40.00n
XX2 net21 B2 VDD VNW PHVT11LL_CKT W=0.26u L=40.00n
XX7 ZN B1 net16 VNW PHVT11LL_CKT W=0.86u L=40.00n
XX1 ZN A VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
XX0 net16 net21 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
.ENDS OAI2XB1V3_12TH40
.SUBCKT OAI2XB1V4_12TH40 A B1 B2 ZN VDD VSS
XX3 net21 B2 VSS VPW NHVT11LL_CKT W=0.305u L=40.00n
XX6 net29 net21 VSS VPW NHVT11LL_CKT W=1.01u L=40.00n
XX5 net29 B1 VSS VPW NHVT11LL_CKT W=1.01u L=40.00n
XX8 ZN A net29 VPW NHVT11LL_CKT W=1.01u L=40.00n
XX2 net21 B2 VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX7 ZN B1 net16 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 ZN A VDD VNW PHVT11LL_CKT W=0.65u L=40.00n
XX0 net16 net21 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS OAI2XB1V4_12TH40
.SUBCKT OAI2XB1V6_12TH40 A B1 B2 ZN VDD VSS
XX3 net21 B2 VSS VPW NHVT11LL_CKT W=0.44u L=40.00n
XX6 net29 net21 VSS VPW NHVT11LL_CKT W=1.515u L=40.00n
XX5 net29 B1 VSS VPW NHVT11LL_CKT W=1.515u L=40.00n
XX8 ZN A net29 VPW NHVT11LL_CKT W=1.515u L=40.00n
XX2 net21 B2 VDD VNW PHVT11LL_CKT W=0.505u L=40.00n
XX7 ZN B1 net16 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX1 ZN A VDD VNW PHVT11LL_CKT W=0.98u L=40.00n
XX0 net16 net21 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS OAI2XB1V6_12TH40
.SUBCKT OAI2XB1V8_12TH40 A B1 B2 ZN VDD VSS
XX3 net21 B2 VSS VPW NHVT11LL_CKT W=0.59u L=40.00n
XX6 net29 net21 VSS VPW NHVT11LL_CKT W=2.02u L=40.00n
XX5 net29 B1 VSS VPW NHVT11LL_CKT W=2.02u L=40.00n
XX8 ZN A net29 VPW NHVT11LL_CKT W=2.02u L=40.00n
XX2 net21 B2 VDD VNW PHVT11LL_CKT W=0.67u L=40.00n
XX7 ZN B1 net16 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 ZN A VDD VNW PHVT11LL_CKT W=1.3u L=40.00n
XX0 net16 net21 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS OAI2XB1V8_12TH40
.SUBCKT OAI31V0_12TH40 A1 A2 A3 B ZN VDD VSS
XX2 net6 A3 VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX5 net6 A1 VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX6 net6 A2 VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX8 ZN B net6 VPW NHVT11LL_CKT W=0.185u L=40.00n
XX3 net29 A3 VDD VNW PHVT11LL_CKT W=0.325u L=40.00n
XX0 net33 A2 net29 VNW PHVT11LL_CKT W=0.325u L=40.00n
XX7 ZN A1 net33 VNW PHVT11LL_CKT W=0.325u L=40.00n
XX1 ZN B VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
.ENDS OAI31V0_12TH40
.SUBCKT OAI31V12_12TH40 A1 A2 A3 B ZN VDD VSS
XX2 net6 A3 VSS VPW NHVT11LL_CKT W=2.1u L=40.00n
XX5 net6 A1 VSS VPW NHVT11LL_CKT W=2.1u L=40.00n
XX6 net6 A2 VSS VPW NHVT11LL_CKT W=2.1u L=40.00n
XX8 ZN B net6 VPW NHVT11LL_CKT W=2.1u L=40.00n
XX3 net29 A3 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX0 net33 A2 net29 VNW PHVT11LL_CKT W=3.66u L=40.00n
XX7 ZN A1 net33 VNW PHVT11LL_CKT W=3.66u L=40.00n
XX1 ZN B VDD VNW PHVT11LL_CKT W=1.35u L=40.00n
.ENDS OAI31V12_12TH40
.SUBCKT OAI31V1_12TH40 A1 A2 A3 B ZN VDD VSS
XX2 net6 A3 VSS VPW NHVT11LL_CKT W=0.245u L=40.00n
XX5 net6 A1 VSS VPW NHVT11LL_CKT W=0.245u L=40.00n
XX6 net6 A2 VSS VPW NHVT11LL_CKT W=0.245u L=40.00n
XX8 ZN B net6 VPW NHVT11LL_CKT W=0.245u L=40.00n
XX3 net29 A3 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX0 net33 A2 net29 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX7 ZN A1 net33 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX1 ZN B VDD VNW PHVT11LL_CKT W=0.16u L=40.00n
.ENDS OAI31V1_12TH40
.SUBCKT OAI31V2_12TH40 A1 A2 A3 B ZN VDD VSS
XX2 net6 A3 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX5 net6 A1 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX6 net6 A2 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX8 ZN B net6 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX3 net29 A3 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX0 net33 A2 net29 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX7 ZN A1 net33 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 ZN B VDD VNW PHVT11LL_CKT W=225.00n L=40.00n
.ENDS OAI31V2_12TH40
.SUBCKT OAI31V3_12TH40 A1 A2 A3 B ZN VDD VSS
XX2 net6 A3 VSS VPW NHVT11LL_CKT W=0.49u L=40.00n
XX5 net6 A1 VSS VPW NHVT11LL_CKT W=0.49u L=40.00n
XX6 net6 A2 VSS VPW NHVT11LL_CKT W=0.49u L=40.00n
XX8 ZN B net6 VPW NHVT11LL_CKT W=0.49u L=40.00n
XX3 net29 A3 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX0 net33 A2 net29 VNW PHVT11LL_CKT W=0.86u L=40.00n
XX7 ZN A1 net33 VNW PHVT11LL_CKT W=0.86u L=40.00n
XX1 ZN B VDD VNW PHVT11LL_CKT W=0.32u L=40.00n
.ENDS OAI31V3_12TH40
.SUBCKT OAI31V4_12TH40 A1 A2 A3 B ZN VDD VSS
XX2 net6 A3 VSS VPW NHVT11LL_CKT W=0.7u L=40.00n
XX5 net6 A1 VSS VPW NHVT11LL_CKT W=0.7u L=40.00n
XX6 net6 A2 VSS VPW NHVT11LL_CKT W=0.7u L=40.00n
XX8 ZN B net6 VPW NHVT11LL_CKT W=0.7u L=40.00n
XX3 net29 A3 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 net33 A2 net29 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX7 ZN A1 net33 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 ZN B VDD VNW PHVT11LL_CKT W=0.45u L=40.00n
.ENDS OAI31V4_12TH40
.SUBCKT OAI31V6_12TH40 A1 A2 A3 B ZN VDD VSS
XX2 net6 A3 VSS VPW NHVT11LL_CKT W=1.05u L=40.00n
XX5 net6 A1 VSS VPW NHVT11LL_CKT W=1.05u L=40.00n
XX6 net6 A2 VSS VPW NHVT11LL_CKT W=1.05u L=40.00n
XX8 ZN B net6 VPW NHVT11LL_CKT W=1.05u L=40.00n
XX3 net29 A3 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX0 net33 A2 net29 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX7 ZN A1 net33 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX1 ZN B VDD VNW PHVT11LL_CKT W=0.68u L=40.00n
.ENDS OAI31V6_12TH40
.SUBCKT OAI31V8_12TH40 A1 A2 A3 B ZN VDD VSS
XX2 net6 A3 VSS VPW NHVT11LL_CKT W=1.4u L=40.00n
XX5 net6 A1 VSS VPW NHVT11LL_CKT W=1.4u L=40.00n
XX6 net6 A2 VSS VPW NHVT11LL_CKT W=1.4u L=40.00n
XX8 ZN B net6 VPW NHVT11LL_CKT W=1.4u L=40.00n
XX3 net29 A3 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX0 net33 A2 net29 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX7 ZN A1 net33 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 ZN B VDD VNW PHVT11LL_CKT W=0.9u L=40.00n
.ENDS OAI31V8_12TH40
.SUBCKT OAI32V1_12TH40 A1 A2 A3 B1 B2 ZN VDD VSS
XX9 ZN B2 net6 VPW NHVT11LL_CKT W=250.00n L=40.00n
XX2 net6 A3 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX5 net6 A1 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX6 net6 A2 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX8 ZN B1 net6 VPW NHVT11LL_CKT W=250.00n L=40.00n
XX4 net055 B2 VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
XX3 net29 A3 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX0 net33 A2 net29 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX7 ZN A1 net33 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX1 ZN B1 net055 VNW PHVT11LL_CKT W=310.00n L=40.00n
.ENDS OAI32V1_12TH40
.SUBCKT OAI32V2_12TH40 A1 A2 A3 B1 B2 ZN VDD VSS
XX9 ZN B2 net6 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX2 net6 A3 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX5 net6 A1 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX6 net6 A2 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX8 ZN B1 net6 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX4 net055 B2 VDD VNW PHVT11LL_CKT W=460.00n L=40.00n
XX3 net29 A3 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX0 net33 A2 net29 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX7 ZN A1 net33 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 ZN B1 net055 VNW PHVT11LL_CKT W=460.00n L=40.00n
.ENDS OAI32V2_12TH40
.SUBCKT OAI32V4_12TH40 A1 A2 A3 B1 B2 ZN VDD VSS
XX9 ZN B2 net6 VPW NHVT11LL_CKT W=700.00n L=40.00n
XX2 net6 A3 VSS VPW NHVT11LL_CKT W=700.00n L=40.00n
XX5 net6 A1 VSS VPW NHVT11LL_CKT W=700.00n L=40.00n
XX6 net6 A2 VSS VPW NHVT11LL_CKT W=700.00n L=40.00n
XX8 ZN B1 net6 VPW NHVT11LL_CKT W=700.00n L=40.00n
XX4 net055 B2 VDD VNW PHVT11LL_CKT W=920.00n L=40.00n
XX3 net29 A3 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 net33 A2 net29 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX7 ZN A1 net33 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 ZN B1 net055 VNW PHVT11LL_CKT W=920.00n L=40.00n
.ENDS OAI32V4_12TH40
.SUBCKT OAI32V8_12TH40 A1 A2 A3 B1 B2 ZN VDD VSS
XX9 ZN B2 net6 VPW NHVT11LL_CKT W=1.4u L=40.00n
XX2 net6 A3 VSS VPW NHVT11LL_CKT W=1.4u L=40.00n
XX5 net6 A1 VSS VPW NHVT11LL_CKT W=1.4u L=40.00n
XX6 net6 A2 VSS VPW NHVT11LL_CKT W=1.4u L=40.00n
XX8 ZN B1 net6 VPW NHVT11LL_CKT W=1.4u L=40.00n
XX4 net055 B2 VDD VNW PHVT11LL_CKT W=1.84u L=40.00n
XX3 net29 A3 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX0 net33 A2 net29 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX7 ZN A1 net33 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 ZN B1 net055 VNW PHVT11LL_CKT W=1.84u L=40.00n
.ENDS OAI32V8_12TH40
.SUBCKT OAI33V1_12TH40 A1 A2 A3 B1 B2 B3 ZN VDD VSS
XX11 ZN B3 net6 VPW NHVT11LL_CKT W=250.00n L=40.00n
XX9 ZN B2 net6 VPW NHVT11LL_CKT W=250.00n L=40.00n
XX2 net6 A3 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX5 net6 A1 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX6 net6 A2 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX8 ZN B1 net6 VPW NHVT11LL_CKT W=250.00n L=40.00n
XX10 net050 B3 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX4 net055 B2 net050 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX3 net29 A3 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX0 net33 A2 net29 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX7 ZN A1 net33 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX1 ZN B1 net055 VNW PHVT11LL_CKT W=430.00n L=40.00n
.ENDS OAI33V1_12TH40
.SUBCKT OAI33V2_12TH40 A1 A2 A3 B1 B2 B3 ZN VDD VSS
XX11 ZN B3 net6 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX9 ZN B2 net6 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX2 net6 A3 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX5 net6 A1 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX6 net6 A2 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX8 ZN B1 net6 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX10 net050 B3 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX4 net055 B2 net050 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX3 net29 A3 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX0 net33 A2 net29 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX7 ZN A1 net33 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 ZN B1 net055 VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS OAI33V2_12TH40
.SUBCKT OAI33V4_12TH40 A1 A2 A3 B1 B2 B3 ZN VDD VSS
XX11 ZN B3 net6 VPW NHVT11LL_CKT W=700.00n L=40.00n
XX9 ZN B2 net6 VPW NHVT11LL_CKT W=700.00n L=40.00n
XX2 net6 A3 VSS VPW NHVT11LL_CKT W=700.00n L=40.00n
XX5 net6 A1 VSS VPW NHVT11LL_CKT W=700.00n L=40.00n
XX6 net6 A2 VSS VPW NHVT11LL_CKT W=700.00n L=40.00n
XX8 ZN B1 net6 VPW NHVT11LL_CKT W=700.00n L=40.00n
XX10 net050 B3 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX4 net055 B2 net050 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX3 net29 A3 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 net33 A2 net29 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX7 ZN A1 net33 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 ZN B1 net055 VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS OAI33V4_12TH40
.SUBCKT OAI33V8_12TH40 A1 A2 A3 B1 B2 B3 ZN VDD VSS
XX11 ZN B3 net6 VPW NHVT11LL_CKT W=1.4u L=40.00n
XX9 ZN B2 net6 VPW NHVT11LL_CKT W=1.4u L=40.00n
XX2 net6 A3 VSS VPW NHVT11LL_CKT W=1.4u L=40.00n
XX5 net6 A1 VSS VPW NHVT11LL_CKT W=1.4u L=40.00n
XX6 net6 A2 VSS VPW NHVT11LL_CKT W=1.4u L=40.00n
XX8 ZN B1 net6 VPW NHVT11LL_CKT W=1.4u L=40.00n
XX10 net050 B3 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX4 net055 B2 net050 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX3 net29 A3 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX0 net33 A2 net29 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX7 ZN A1 net33 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 ZN B1 net055 VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS OAI33V8_12TH40
.SUBCKT OAO211V1_12TH40 A1 A2 B C Z VDD VSS
XX6 net031 C VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX2 net10 A1 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX0 net10 A2 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX5 net031 B net10 VPW NHVT11LL_CKT W=250.00n L=40.00n
XX8 Z net031 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX7 Z net031 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX4 net031 C net30 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX3 net33 A2 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX9 net30 A1 net33 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX1 net30 B VDD VNW PHVT11LL_CKT W=330.00n L=40.00n
.ENDS OAO211V1_12TH40
.SUBCKT OAO211V2_12TH40 A1 A2 B C Z VDD VSS
XX6 net031 C VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX2 net10 A1 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX0 net10 A2 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX5 net031 B net10 VPW NHVT11LL_CKT W=350.00n L=40.00n
XX8 Z net031 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX7 Z net031 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX4 net031 C net30 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX3 net33 A2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX9 net30 A1 net33 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 net30 B VDD VNW PHVT11LL_CKT W=450.00n L=40.00n
.ENDS OAO211V2_12TH40
.SUBCKT OAO211V4_12TH40 A1 A2 B C Z VDD VSS
XX6 net031 C VSS VPW NHVT11LL_CKT W=440.00n L=40.00n
XX2 net10 A1 VSS VPW NHVT11LL_CKT W=700.00n L=40.00n
XX0 net10 A2 VSS VPW NHVT11LL_CKT W=700.00n L=40.00n
XX5 net031 B net10 VPW NHVT11LL_CKT W=700.00n L=40.00n
XX8 Z net031 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX7 Z net031 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX4 net031 C net30 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX3 net33 A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX9 net30 A1 net33 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 net30 B VDD VNW PHVT11LL_CKT W=900.00n L=40.00n
.ENDS OAO211V4_12TH40
.SUBCKT OAO211V8_12TH40 A1 A2 B C Z VDD VSS
XX6 net031 C VSS VPW NHVT11LL_CKT W=880.00n L=40.00n
XX2 net10 A1 VSS VPW NHVT11LL_CKT W=1.4u L=40.00n
XX0 net10 A2 VSS VPW NHVT11LL_CKT W=1.4u L=40.00n
XX5 net031 B net10 VPW NHVT11LL_CKT W=1.4u L=40.00n
XX8 Z net031 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX7 Z net031 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX4 net031 C net30 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX3 net33 A2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX9 net30 A1 net33 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 net30 B VDD VNW PHVT11LL_CKT W=1.84u L=40.00n
.ENDS OAO211V8_12TH40
.SUBCKT OAOAI2111V1_12TH40 A1 A2 B C D ZN VDD VSS
XX10 net31 A2 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX9 net31 A1 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX6 net35 B net31 VPW NHVT11LL_CKT W=380.00n L=40.00n
XX8 net35 C VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX5 ZN D net35 VPW NHVT11LL_CKT W=0.375u L=40.00n
XX4 ZN C net11 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX3 net11 A1 net14 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX2 ZN D VDD VNW PHVT11LL_CKT W=220.00n L=40.00n
XX1 net11 B VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
XX0 net14 A2 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
.ENDS OAOAI2111V1_12TH40
.SUBCKT OAOAI2111V2_12TH40 A1 A2 B C D ZN VDD VSS
XX10 net31 A2 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX9 net31 A1 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX6 net35 B net31 VPW NHVT11LL_CKT W=540.00n L=40.00n
XX8 net35 C VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX5 ZN D net35 VPW NHVT11LL_CKT W=540.00n L=40.00n
XX4 ZN C net11 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX3 net11 A1 net14 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX2 ZN D VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
XX1 net11 B VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX0 net14 A2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS OAOAI2111V2_12TH40
.SUBCKT OAOAI2111V4_12TH40 A1 A2 B C D ZN VDD VSS
XX10 net31 A2 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX9 net31 A1 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX6 net35 B net31 VPW NHVT11LL_CKT W=1.08u L=40.00n
XX8 net35 C VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX5 ZN D net35 VPW NHVT11LL_CKT W=1.08u L=40.00n
XX4 ZN C net11 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX3 net11 A1 net14 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX2 ZN D VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 net11 B VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX0 net14 A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS OAOAI2111V4_12TH40
.SUBCKT OAOAI2111V8_12TH40 A1 A2 B C D ZN VDD VSS
XX10 net31 A2 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX9 net31 A1 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX6 net35 B net31 VPW NHVT11LL_CKT W=2.16u L=40.00n
XX8 net35 C VSS VPW NHVT11LL_CKT W=1.52u L=40.00n
XX5 ZN D net35 VPW NHVT11LL_CKT W=2.16u L=40.00n
XX4 ZN C net11 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX3 net11 A1 net14 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX2 ZN D VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 net11 B VDD VNW PHVT11LL_CKT W=1.72u L=40.00n
XX0 net14 A2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS OAOAI2111V8_12TH40
.SUBCKT OAOAOAI211111V1_12TH40 A1 A2 B C D E F ZN VDD VSS
XX13 net29 E VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX12 net25 C VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX11 net21 A2 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX10 net21 A1 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX9 net25 B net21 VPW NHVT11LL_CKT W=380.00n L=40.00n
XX8 net29 D net25 VPW NHVT11LL_CKT W=380.00n L=40.00n
XX7 ZN F net29 VPW NHVT11LL_CKT W=380.00n L=40.00n
XX5 net64 C net53 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX3 net64 D VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
XX2 net53 B VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX4 ZN F VDD VNW PHVT11LL_CKT W=220.00n L=40.00n
XX1 net53 A1 net56 VNW PHVT11LL_CKT W=430.00n L=40.00n
XX0 net56 A2 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX6 ZN E net64 VNW PHVT11LL_CKT W=430.00n L=40.00n
.ENDS OAOAOAI211111V1_12TH40
.SUBCKT OAOAOAI211111V2_12TH40 A1 A2 B C D E F ZN VDD VSS
XX13 net29 E VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX12 net25 C VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX11 net21 A2 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX10 net21 A1 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX9 net25 B net21 VPW NHVT11LL_CKT W=540.00n L=40.00n
XX8 net29 D net25 VPW NHVT11LL_CKT W=540.00n L=40.00n
XX7 ZN F net29 VPW NHVT11LL_CKT W=540.00n L=40.00n
XX5 net64 C net53 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX3 net64 D VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX2 net53 B VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX4 ZN F VDD VNW PHVT11LL_CKT W=310.00n L=40.00n
XX1 net53 A1 net56 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX0 net56 A2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX6 ZN E net64 VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS OAOAOAI211111V2_12TH40
.SUBCKT OAOAOAI211111V4_12TH40 A1 A2 B C D E F ZN VDD VSS
XX13 net29 E VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX12 net25 C VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX11 net21 A2 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX10 net21 A1 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX9 net25 B net21 VPW NHVT11LL_CKT W=1.08u L=40.00n
XX8 net29 D net25 VPW NHVT11LL_CKT W=1.08u L=40.00n
XX7 ZN F net29 VPW NHVT11LL_CKT W=1.08u L=40.00n
XX5 net64 C net53 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX3 net64 D VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX2 net53 B VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX4 ZN F VDD VNW PHVT11LL_CKT W=620.00n L=40.00n
XX1 net53 A1 net56 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 net56 A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX6 ZN E net64 VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS OAOAOAI211111V4_12TH40
.SUBCKT OAOAOAI211111V8_12TH40 A1 A2 B C D E F ZN VDD VSS
XX13 net29 E VSS VPW NHVT11LL_CKT W=1.52u L=40.00n
XX12 net25 C VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX11 net21 A2 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX10 net21 A1 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX9 net25 B net21 VPW NHVT11LL_CKT W=2.16u L=40.00n
XX8 net29 D net25 VPW NHVT11LL_CKT W=2.16u L=40.00n
XX7 ZN F net29 VPW NHVT11LL_CKT W=2.16u L=40.00n
XX5 net64 C net53 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX3 net64 D VDD VNW PHVT11LL_CKT W=1.72u L=40.00n
XX2 net53 B VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX4 ZN F VDD VNW PHVT11LL_CKT W=1.24u L=40.00n
XX1 net53 A1 net56 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX0 net56 A2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX6 ZN E net64 VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS OAOAOAI211111V8_12TH40
.SUBCKT OAOI211V0_12TH40 A1 A2 B C ZN VDD VSS
XX6 ZN C VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX2 net10 A1 VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX0 net10 A2 VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX5 ZN B net10 VPW NHVT11LL_CKT W=0.21u L=40.00n
XX4 ZN C net30 VNW PHVT11LL_CKT W=0.365u L=40.00n
XX3 net33 A2 VDD VNW PHVT11LL_CKT W=0.365u L=40.00n
XX9 net30 A1 net33 VNW PHVT11LL_CKT W=0.365u L=40.00n
XX1 net30 B VDD VNW PHVT11LL_CKT W=0.255u L=40.00n
.ENDS OAOI211V0_12TH40
.SUBCKT OAOI211V12_12TH40 A1 A2 B C ZN VDD VSS
XX6 ZN C VSS VPW NHVT11LL_CKT W=1.2u L=40.00n
XX2 net10 A1 VSS VPW NHVT11LL_CKT W=2.1u L=40.00n
XX0 net10 A2 VSS VPW NHVT11LL_CKT W=2.1u L=40.00n
XX5 ZN B net10 VPW NHVT11LL_CKT W=2.1u L=40.00n
XX4 ZN C net30 VNW PHVT11LL_CKT W=3.66u L=40.00n
XX3 net33 A2 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
XX9 net30 A1 net33 VNW PHVT11LL_CKT W=3.66u L=40.00n
XX1 net30 B VDD VNW PHVT11LL_CKT W=2.55u L=40.00n
.ENDS OAOI211V12_12TH40
.SUBCKT OAOI211V1_12TH40 A1 A2 B C ZN VDD VSS
XX6 ZN C VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX2 net10 A1 VSS VPW NHVT11LL_CKT W=0.245u L=40.00n
XX0 net10 A2 VSS VPW NHVT11LL_CKT W=0.245u L=40.00n
XX5 ZN B net10 VPW NHVT11LL_CKT W=0.245u L=40.00n
XX4 ZN C net30 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX3 net33 A2 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX9 net30 A1 net33 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX1 net30 B VDD VNW PHVT11LL_CKT W=0.3u L=40.00n
.ENDS OAOI211V1_12TH40
.SUBCKT OAOI211V2_12TH40 A1 A2 B C ZN VDD VSS
XX6 ZN C VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX2 net10 A1 VSS VPW NHVT11LL_CKT W=0.355u L=40.00n
XX0 net10 A2 VSS VPW NHVT11LL_CKT W=0.355u L=40.00n
XX5 ZN B net10 VPW NHVT11LL_CKT W=0.355u L=40.00n
XX4 ZN C net30 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX3 net33 A2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX9 net30 A1 net33 VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 net30 B VDD VNW PHVT11LL_CKT W=425.00n L=40.00n
.ENDS OAOI211V2_12TH40
.SUBCKT OAOI211V3_12TH40 A1 A2 B C ZN VDD VSS
XX6 ZN C VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX2 net10 A1 VSS VPW NHVT11LL_CKT W=0.49u L=40.00n
XX0 net10 A2 VSS VPW NHVT11LL_CKT W=0.49u L=40.00n
XX5 ZN B net10 VPW NHVT11LL_CKT W=0.49u L=40.00n
XX4 ZN C net30 VNW PHVT11LL_CKT W=0.86u L=40.00n
XX3 net33 A2 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX9 net30 A1 net33 VNW PHVT11LL_CKT W=0.86u L=40.00n
XX1 net30 B VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
.ENDS OAOI211V3_12TH40
.SUBCKT OAOI211V4_12TH40 A1 A2 B C ZN VDD VSS
XX6 ZN C VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX2 net10 A1 VSS VPW NHVT11LL_CKT W=0.7u L=40.00n
XX0 net10 A2 VSS VPW NHVT11LL_CKT W=0.7u L=40.00n
XX5 ZN B net10 VPW NHVT11LL_CKT W=0.7u L=40.00n
XX4 ZN C net30 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX3 net33 A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX9 net30 A1 net33 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 net30 B VDD VNW PHVT11LL_CKT W=0.85u L=40.00n
.ENDS OAOI211V4_12TH40
.SUBCKT OAOI211V6_12TH40 A1 A2 B C ZN VDD VSS
XX6 ZN C VSS VPW NHVT11LL_CKT W=0.6u L=40.00n
XX2 net10 A1 VSS VPW NHVT11LL_CKT W=1.05u L=40.00n
XX0 net10 A2 VSS VPW NHVT11LL_CKT W=1.05u L=40.00n
XX5 ZN B net10 VPW NHVT11LL_CKT W=1.05u L=40.00n
XX4 ZN C net30 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX3 net33 A2 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX9 net30 A1 net33 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX1 net30 B VDD VNW PHVT11LL_CKT W=1.275u L=40.00n
.ENDS OAOI211V6_12TH40
.SUBCKT OAOI211V8_12TH40 A1 A2 B C ZN VDD VSS
XX6 ZN C VSS VPW NHVT11LL_CKT W=0.8u L=40.00n
XX2 net10 A1 VSS VPW NHVT11LL_CKT W=1.4u L=40.00n
XX0 net10 A2 VSS VPW NHVT11LL_CKT W=1.4u L=40.00n
XX5 ZN B net10 VPW NHVT11LL_CKT W=1.4u L=40.00n
XX4 ZN C net30 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX3 net33 A2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX9 net30 A1 net33 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 net30 B VDD VNW PHVT11LL_CKT W=1.7u L=40.00n
.ENDS OAOI211V8_12TH40
.SUBCKT OR2V0_12TH40 A1 A2 Z VDD VSS
XX5 net8 A1 VSS VPW NHVT11LL_CKT W=0.125u L=40.00n
XX6 net8 A2 VSS VPW NHVT11LL_CKT W=0.125u L=40.00n
XX8 Z net8 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX0 net23 A2 VDD VNW PHVT11LL_CKT W=0.27u L=40.00n
XX7 net8 A1 net23 VNW PHVT11LL_CKT W=0.27u L=40.00n
XX1 Z net8 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
.ENDS OR2V0_12TH40
.SUBCKT OR2V10RD_12TH40 A1 A2 Z VDD VSS
XX5 net8 A1 VSS VPW NHVT11LL_CKT W=1.82u L=40.00n
XX6 net8 A2 VSS VPW NHVT11LL_CKT W=1.82u L=40.00n
XX8 Z net8 VSS VPW NHVT11LL_CKT W=2.7u L=40.00n
XX0 net23 A2 VDD VNW PHVT11LL_CKT W=5.49u L=40.00n
XX7 net8 A1 net23 VNW PHVT11LL_CKT W=5.49u L=40.00n
XX1 Z net8 VDD VNW PHVT11LL_CKT W=3.05u L=40.00n
.ENDS OR2V10RD_12TH40
.SUBCKT OR2V12_12TH40 A1 A2 Z VDD VSS
XX5 net8 A1 VSS VPW NHVT11LL_CKT W=1.12u L=40.00n
XX6 net8 A2 VSS VPW NHVT11LL_CKT W=1.12u L=40.00n
XX8 Z net8 VSS VPW NHVT11LL_CKT W=3.21u L=40.00n
XX0 net23 A2 VDD VNW PHVT11LL_CKT W=2.4u L=40.00n
XX7 net8 A1 net23 VNW PHVT11LL_CKT W=2.4u L=40.00n
XX1 Z net8 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
.ENDS OR2V12_12TH40
.SUBCKT OR2V16_12TH40 A1 A2 Z VDD VSS
XX5 net8 A1 VSS VPW NHVT11LL_CKT W=1.53u L=40.00n
XX6 net8 A2 VSS VPW NHVT11LL_CKT W=1.53u L=40.00n
XX8 Z net8 VSS VPW NHVT11LL_CKT W=4.28u L=40.00n
XX0 net23 A2 VDD VNW PHVT11LL_CKT W=3.27u L=40.00n
XX7 net8 A1 net23 VNW PHVT11LL_CKT W=3.27u L=40.00n
XX1 Z net8 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
.ENDS OR2V16_12TH40
.SUBCKT OR2V1RD_12TH40 A1 A2 Z VDD VSS
XX5 net8 A1 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX6 net8 A2 VSS VPW NHVT11LL_CKT W=250.00n L=40.00n
XX8 Z net8 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX0 net23 A2 VDD VNW PHVT11LL_CKT W=760.00n L=40.00n
XX7 net8 A1 net23 VNW PHVT11LL_CKT W=760.00n L=40.00n
XX1 Z net8 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
.ENDS OR2V1RD_12TH40
.SUBCKT OR2V1_12TH40 A1 A2 Z VDD VSS
XX5 net8 A1 VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX6 net8 A2 VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX8 Z net8 VSS VPW NHVT11LL_CKT W=0.375u L=40.00n
XX0 net23 A2 VDD VNW PHVT11LL_CKT W=0.34u L=40.00n
XX7 net8 A1 net23 VNW PHVT11LL_CKT W=0.34u L=40.00n
XX1 Z net8 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
.ENDS OR2V1_12TH40
.SUBCKT OR2V22_12TH40 A1 A2 Z VDD VSS
XX5 net8 A1 VSS VPW NHVT11LL_CKT W=1.995u L=40.00n
XX6 net8 A2 VSS VPW NHVT11LL_CKT W=1.995u L=40.00n
XX8 Z net8 VSS VPW NHVT11LL_CKT W=5.885u L=40.00n
XX0 net23 A2 VDD VNW PHVT11LL_CKT W=4.27u L=40.00n
XX7 net8 A1 net23 VNW PHVT11LL_CKT W=4.27u L=40.00n
XX1 Z net8 VDD VNW PHVT11LL_CKT W=6.71u L=40.00n
.ENDS OR2V22_12TH40
.SUBCKT OR2V2RD_12TH40 A1 A2 Z VDD VSS
XX5 net8 A1 VSS VPW NHVT11LL_CKT W=360.00n L=40.00n
XX6 net8 A2 VSS VPW NHVT11LL_CKT W=360.00n L=40.00n
XX8 Z net8 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX0 net23 A2 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX7 net8 A1 net23 VNW PHVT11LL_CKT W=1.08u L=40.00n
XX1 Z net8 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS OR2V2RD_12TH40
.SUBCKT OR2V2_12TH40 A1 A2 Z VDD VSS
XX5 net8 A1 VSS VPW NHVT11LL_CKT W=205.00n L=40.00n
XX6 net8 A2 VSS VPW NHVT11LL_CKT W=205.00n L=40.00n
XX8 Z net8 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX0 net23 A2 VDD VNW PHVT11LL_CKT W=435.00n L=40.00n
XX7 net8 A1 net23 VNW PHVT11LL_CKT W=435.00n L=40.00n
XX1 Z net8 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS OR2V2_12TH40
.SUBCKT OR2V3_12TH40 A1 A2 Z VDD VSS
XX5 net8 A1 VSS VPW NHVT11LL_CKT W=275.00n L=40.00n
XX6 net8 A2 VSS VPW NHVT11LL_CKT W=275.00n L=40.00n
XX8 Z net8 VSS VPW NHVT11LL_CKT W=760.00n L=40.00n
XX0 net23 A2 VDD VNW PHVT11LL_CKT W=580.00n L=40.00n
XX7 net8 A1 net23 VNW PHVT11LL_CKT W=580.00n L=40.00n
XX1 Z net8 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
.ENDS OR2V3_12TH40
.SUBCKT OR2V4RD_12TH40 A1 A2 Z VDD VSS
XX5 net8 A1 VSS VPW NHVT11LL_CKT W=720.00n L=40.00n
XX6 net8 A2 VSS VPW NHVT11LL_CKT W=720.00n L=40.00n
XX8 Z net8 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX0 net23 A2 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
XX7 net8 A1 net23 VNW PHVT11LL_CKT W=2.16u L=40.00n
XX1 Z net8 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS OR2V4RD_12TH40
.SUBCKT OR2V4_12TH40 A1 A2 Z VDD VSS
XX5 net8 A1 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX6 net8 A2 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX8 Z net8 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX0 net23 A2 VDD VNW PHVT11LL_CKT W=0.84u L=40.00n
XX7 net8 A1 net23 VNW PHVT11LL_CKT W=0.84u L=40.00n
XX1 Z net8 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS OR2V4_12TH40
.SUBCKT OR2V6RD_12TH40 A1 A2 Z VDD VSS
XX5 net8 A1 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX6 net8 A2 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX8 Z net8 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX0 net23 A2 VDD VNW PHVT11LL_CKT W=3.24u L=40.00n
XX7 net8 A1 net23 VNW PHVT11LL_CKT W=3.24u L=40.00n
XX1 Z net8 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS OR2V6RD_12TH40
.SUBCKT OR2V6_12TH40 A1 A2 Z VDD VSS
XX5 net8 A1 VSS VPW NHVT11LL_CKT W=0.56u L=40.00n
XX6 net8 A2 VSS VPW NHVT11LL_CKT W=0.56u L=40.00n
XX8 Z net8 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX0 net23 A2 VDD VNW PHVT11LL_CKT W=1.19u L=40.00n
XX7 net8 A1 net23 VNW PHVT11LL_CKT W=1.19u L=40.00n
XX1 Z net8 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS OR2V6_12TH40
.SUBCKT OR2V8RD_12TH40 A1 A2 Z VDD VSS
XX5 net8 A1 VSS VPW NHVT11LL_CKT W=1.42u L=40.00n
XX6 net8 A2 VSS VPW NHVT11LL_CKT W=1.42u L=40.00n
XX8 Z net8 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX0 net23 A2 VDD VNW PHVT11LL_CKT W=4.27u L=40.00n
XX7 net8 A1 net23 VNW PHVT11LL_CKT W=4.27u L=40.00n
XX1 Z net8 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS OR2V8RD_12TH40
.SUBCKT OR2V8_12TH40 A1 A2 Z VDD VSS
XX5 net8 A1 VSS VPW NHVT11LL_CKT W=0.765u L=40.00n
XX6 net8 A2 VSS VPW NHVT11LL_CKT W=0.765u L=40.00n
XX8 Z net8 VSS VPW NHVT11LL_CKT W=2.14u L=40.00n
XX0 net23 A2 VDD VNW PHVT11LL_CKT W=1.62u L=40.00n
XX7 net8 A1 net23 VNW PHVT11LL_CKT W=1.62u L=40.00n
XX1 Z net8 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS OR2V8_12TH40
.SUBCKT OR3V0_12TH40 A1 A2 A3 Z VDD VSS
XX3 net8 A3 VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX5 net8 A1 VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX6 net8 A2 VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX8 Z net8 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX2 net064 A3 VDD VNW PHVT11LL_CKT W=0.505u L=40.00n
XX0 net23 A2 net064 VNW PHVT11LL_CKT W=0.505u L=40.00n
XX7 net8 A1 net23 VNW PHVT11LL_CKT W=0.505u L=40.00n
XX1 Z net8 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
.ENDS OR3V0_12TH40
.SUBCKT OR3V10RD_12TH40 A1 A2 A3 Z VDD VSS
XX1 Z A3N VDD VNW PHVT11LL_CKT W=2.7u L=40.00n
XX0 net48 A1 net23 VNW PHVT11LL_CKT W=5.4u L=40.00n
XX4 net23 A2 VDD VNW PHVT11LL_CKT W=5.4u L=40.00n
XX8 A3N A3 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX3 Z net48 VDD VNW PHVT11LL_CKT W=2.7u L=40.00n
XX9 A3N A3 VSS VPW NHVT11LL_CKT W=1.23u L=40.00n
XX5 net48 A2 VSS VPW NHVT11LL_CKT W=2.00u L=40.00n
XX7 Z net48 net40 VPW NHVT11LL_CKT W=3.05u L=40.00n
XX6 net40 A3N VSS VPW NHVT11LL_CKT W=3.05u L=40.00n
XX2 net48 A1 VSS VPW NHVT11LL_CKT W=2.00u L=40.00n
.ENDS OR3V10RD_12TH40
.SUBCKT OR3V12_12TH40 A1 A2 A3 Z VDD VSS
XX3 net8 A3 VSS VPW NHVT11LL_CKT W=1.44u L=40.00n
XX5 net8 A1 VSS VPW NHVT11LL_CKT W=1.44u L=40.00n
XX6 net8 A2 VSS VPW NHVT11LL_CKT W=1.44u L=40.00n
XX8 Z net8 VSS VPW NHVT11LL_CKT W=3.21u L=40.00n
XX2 net064 A3 VDD VNW PHVT11LL_CKT W=4.64u L=40.00n
XX0 net23 A2 net064 VNW PHVT11LL_CKT W=4.64u L=40.00n
XX7 net8 A1 net23 VNW PHVT11LL_CKT W=4.64u L=40.00n
XX1 Z net8 VDD VNW PHVT11LL_CKT W=3.66u L=40.00n
.ENDS OR3V12_12TH40
.SUBCKT OR3V16_12TH40 A1 A2 A3 Z VDD VSS
XX3 net8 A3 VSS VPW NHVT11LL_CKT W=1.9u L=40.00n
XX5 net8 A1 VSS VPW NHVT11LL_CKT W=1.9u L=40.00n
XX6 net8 A2 VSS VPW NHVT11LL_CKT W=1.9u L=40.00n
XX8 Z net8 VSS VPW NHVT11LL_CKT W=4.28u L=40.00n
XX2 net064 A3 VDD VNW PHVT11LL_CKT W=6.1u L=40.00n
XX0 net23 A2 net064 VNW PHVT11LL_CKT W=6.1u L=40.00n
XX7 net8 A1 net23 VNW PHVT11LL_CKT W=6.1u L=40.00n
XX1 Z net8 VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
.ENDS OR3V16_12TH40
.SUBCKT OR3V1RD_12TH40 A1 A2 A3 Z VDD VSS
XX1 Z A3N VDD VNW PHVT11LL_CKT W=380.00n L=40.00n
XX0 net48 A1 net23 VNW PHVT11LL_CKT W=760.00n L=40.00n
XX4 net23 A2 VDD VNW PHVT11LL_CKT W=760.00n L=40.00n
XX8 A3N A3 VDD VNW PHVT11LL_CKT W=290.00n L=40.00n
XX3 Z net48 VDD VNW PHVT11LL_CKT W=380.00n L=40.00n
XX9 A3N A3 VSS VPW NHVT11LL_CKT W=200.00n L=40.00n
XX5 net48 A2 VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX7 Z net48 net40 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX6 net40 A3N VSS VPW NHVT11LL_CKT W=430.00n L=40.00n
XX2 net48 A1 VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
.ENDS OR3V1RD_12TH40
.SUBCKT OR3V1_12TH40 A1 A2 A3 Z VDD VSS
XX3 net8 A3 VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX5 net8 A1 VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX6 net8 A2 VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX8 Z net8 VSS VPW NHVT11LL_CKT W=0.375u L=40.00n
XX2 net064 A3 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net23 A2 net064 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX7 net8 A1 net23 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX1 Z net8 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
.ENDS OR3V1_12TH40
.SUBCKT OR3V2RD_12TH40 A1 A2 A3 Z VDD VSS
XX1 Z A3N VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX0 net48 A1 net23 VNW PHVT11LL_CKT W=1.08u L=40.00n
XX4 net23 A2 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX8 A3N A3 VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX3 Z net48 VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX9 A3N A3 VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX5 net48 A2 VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX7 Z net48 net40 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX6 net40 A3N VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX2 net48 A1 VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
.ENDS OR3V2RD_12TH40
.SUBCKT OR3V2_12TH40 A1 A2 A3 Z VDD VSS
XX3 net8 A3 VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX5 net8 A1 VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX6 net8 A2 VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX8 Z net8 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX2 net064 A3 VDD VNW PHVT11LL_CKT W=860.00n L=40.00n
XX0 net23 A2 net064 VNW PHVT11LL_CKT W=860.00n L=40.00n
XX7 net8 A1 net23 VNW PHVT11LL_CKT W=860.00n L=40.00n
XX1 Z net8 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS OR3V2_12TH40
.SUBCKT OR3V3_12TH40 A1 A2 A3 Z VDD VSS
XX3 net8 A3 VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX5 net8 A1 VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX6 net8 A2 VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX8 Z net8 VSS VPW NHVT11LL_CKT W=0.75u L=40.00n
XX2 net064 A3 VDD VNW PHVT11LL_CKT W=1.11u L=40.00n
XX0 net23 A2 net064 VNW PHVT11LL_CKT W=1.11u L=40.00n
XX7 net8 A1 net23 VNW PHVT11LL_CKT W=1.11u L=40.00n
XX1 Z net8 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
.ENDS OR3V3_12TH40
.SUBCKT OR3V4RD_12TH40 A1 A2 A3 Z VDD VSS
XX1 Z A3N VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX0 net48 A1 net23 VNW PHVT11LL_CKT W=2.16u L=40.00n
XX4 net23 A2 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
XX8 A3N A3 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX3 Z net48 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX9 A3N A3 VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX5 net48 A2 VSS VPW NHVT11LL_CKT W=800.00n L=40.00n
XX7 Z net48 net40 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX6 net40 A3N VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX2 net48 A1 VSS VPW NHVT11LL_CKT W=800.00n L=40.00n
.ENDS OR3V4RD_12TH40
.SUBCKT OR3V4_12TH40 A1 A2 A3 Z VDD VSS
XX3 net8 A3 VSS VPW NHVT11LL_CKT W=0.48u L=40.00n
XX5 net8 A1 VSS VPW NHVT11LL_CKT W=0.48u L=40.00n
XX6 net8 A2 VSS VPW NHVT11LL_CKT W=0.48u L=40.00n
XX8 Z net8 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX2 net064 A3 VDD VNW PHVT11LL_CKT W=1.53u L=40.00n
XX0 net23 A2 net064 VNW PHVT11LL_CKT W=1.53u L=40.00n
XX7 net8 A1 net23 VNW PHVT11LL_CKT W=1.53u L=40.00n
XX1 Z net8 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS OR3V4_12TH40
.SUBCKT OR3V6RD_12TH40 A1 A2 A3 Z VDD VSS
XX1 Z A3N VDD VNW PHVT11LL_CKT W=1.62u L=40.00n
XX0 net48 A1 net23 VNW PHVT11LL_CKT W=3.24u L=40.00n
XX4 net23 A2 VDD VNW PHVT11LL_CKT W=3.24u L=40.00n
XX8 A3N A3 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX3 Z net48 VDD VNW PHVT11LL_CKT W=1.62u L=40.00n
XX9 A3N A3 VSS VPW NHVT11LL_CKT W=800.00n L=40.00n
XX5 net48 A2 VSS VPW NHVT11LL_CKT W=1.2u L=40.00n
XX7 Z net48 net40 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX6 net40 A3N VSS VPW NHVT11LL_CKT W=1.83u L=40.00n
XX2 net48 A1 VSS VPW NHVT11LL_CKT W=1.2u L=40.00n
.ENDS OR3V6RD_12TH40
.SUBCKT OR3V6_12TH40 A1 A2 A3 Z VDD VSS
XX3 net8 A3 VSS VPW NHVT11LL_CKT W=0.7u L=40.00n
XX5 net8 A1 VSS VPW NHVT11LL_CKT W=0.7u L=40.00n
XX6 net8 A2 VSS VPW NHVT11LL_CKT W=0.7u L=40.00n
XX8 Z net8 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX2 net064 A3 VDD VNW PHVT11LL_CKT W=2.24u L=40.00n
XX0 net23 A2 net064 VNW PHVT11LL_CKT W=2.24u L=40.00n
XX7 net8 A1 net23 VNW PHVT11LL_CKT W=2.24u L=40.00n
XX1 Z net8 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS OR3V6_12TH40
.SUBCKT OR3V8RD_12TH40 A1 A2 A3 Z VDD VSS
XX1 Z A3N VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
XX0 net48 A1 net23 VNW PHVT11LL_CKT W=4.34u L=40.00n
XX4 net23 A2 VDD VNW PHVT11LL_CKT W=4.34u L=40.00n
XX8 A3N A3 VDD VNW PHVT11LL_CKT W=1.59u L=40.00n
XX3 Z net48 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
XX9 A3N A3 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX5 net48 A2 VSS VPW NHVT11LL_CKT W=1.6u L=40.00n
XX7 Z net48 net40 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX6 net40 A3N VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX2 net48 A1 VSS VPW NHVT11LL_CKT W=1.6u L=40.00n
.ENDS OR3V8RD_12TH40
.SUBCKT OR3V8_12TH40 A1 A2 A3 Z VDD VSS
XX3 net8 A3 VSS VPW NHVT11LL_CKT W=0.95u L=40.00n
XX5 net8 A1 VSS VPW NHVT11LL_CKT W=0.95u L=40.00n
XX6 net8 A2 VSS VPW NHVT11LL_CKT W=0.95u L=40.00n
XX8 Z net8 VSS VPW NHVT11LL_CKT W=2.14u L=40.00n
XX2 net064 A3 VDD VNW PHVT11LL_CKT W=3.05u L=40.00n
XX0 net23 A2 net064 VNW PHVT11LL_CKT W=3.05u L=40.00n
XX7 net8 A1 net23 VNW PHVT11LL_CKT W=3.05u L=40.00n
XX1 Z net8 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS OR3V8_12TH40
.SUBCKT OR4V0_12TH40 A1 A2 A3 A4 Z VDD VSS
XX22 DC A4 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX23 DC A3 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX19 Z BA net34 VPW NHVT11LL_CKT W=0.305u L=40.00n
XX6 BA A2 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX5 BA A1 VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX18 net34 DC VSS VPW NHVT11LL_CKT W=0.305u L=40.00n
XX20 DC A3 net21 VNW PHVT11LL_CKT W=0.25u L=40.00n
XX21 net21 A4 VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX16 Z BA VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX17 Z DC VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX0 BA A1 net25 VNW PHVT11LL_CKT W=0.25u L=40.00n
XX2 net25 A2 VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
.ENDS OR4V0_12TH40
.SUBCKT OR4V10RD_12TH40 A1 A2 A3 A4 Z VDD VSS
XX22 DC A4 VSS VPW NHVT11LL_CKT W=2.00u L=40.00n
XX23 DC A3 VSS VPW NHVT11LL_CKT W=2.00u L=40.00n
XX19 Z BA net34 VPW NHVT11LL_CKT W=3.05u L=40.00n
XX6 BA A2 VSS VPW NHVT11LL_CKT W=2.00u L=40.00n
XX5 BA A1 VSS VPW NHVT11LL_CKT W=2.00u L=40.00n
XX18 net34 DC VSS VPW NHVT11LL_CKT W=3.05u L=40.00n
XX20 DC A3 net21 VNW PHVT11LL_CKT W=5.4u L=40.00n
XX21 net21 A4 VDD VNW PHVT11LL_CKT W=5.4u L=40.00n
XX16 Z BA VDD VNW PHVT11LL_CKT W=2.7u L=40.00n
XX17 Z DC VDD VNW PHVT11LL_CKT W=2.7u L=40.00n
XX0 BA A1 net25 VNW PHVT11LL_CKT W=5.4u L=40.00n
XX2 net25 A2 VDD VNW PHVT11LL_CKT W=5.4u L=40.00n
.ENDS OR4V10RD_12TH40
.SUBCKT OR4V12_12TH40 A1 A2 A3 A4 Z VDD VSS
XX22 DC A4 VSS VPW NHVT11LL_CKT W=1.02u L=40.00n
XX23 DC A3 VSS VPW NHVT11LL_CKT W=1.02u L=40.00n
XX19 Z BA net34 VPW NHVT11LL_CKT W=3.66u L=40.00n
XX6 BA A2 VSS VPW NHVT11LL_CKT W=1.02u L=40.00n
XX5 BA A1 VSS VPW NHVT11LL_CKT W=1.02u L=40.00n
XX18 net34 DC VSS VPW NHVT11LL_CKT W=3.66u L=40.00n
XX20 DC A3 net21 VNW PHVT11LL_CKT W=2.16u L=40.00n
XX21 net21 A4 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
XX16 Z BA VDD VNW PHVT11LL_CKT W=2.37u L=40.00n
XX17 Z DC VDD VNW PHVT11LL_CKT W=2.37u L=40.00n
XX0 BA A1 net25 VNW PHVT11LL_CKT W=2.16u L=40.00n
XX2 net25 A2 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
.ENDS OR4V12_12TH40
.SUBCKT OR4V16_12TH40 A1 A2 A3 A4 Z VDD VSS
XX22 DC A4 VSS VPW NHVT11LL_CKT W=1.35u L=40.00n
XX23 DC A3 VSS VPW NHVT11LL_CKT W=1.35u L=40.00n
XX19 Z BA net34 VPW NHVT11LL_CKT W=4.88u L=40.00n
XX6 BA A2 VSS VPW NHVT11LL_CKT W=1.35u L=40.00n
XX5 BA A1 VSS VPW NHVT11LL_CKT W=1.35u L=40.00n
XX18 net34 DC VSS VPW NHVT11LL_CKT W=4.88u L=40.00n
XX20 DC A3 net21 VNW PHVT11LL_CKT W=2.85u L=40.00n
XX21 net21 A4 VDD VNW PHVT11LL_CKT W=2.85u L=40.00n
XX16 Z BA VDD VNW PHVT11LL_CKT W=3.16u L=40.00n
XX17 Z DC VDD VNW PHVT11LL_CKT W=3.16u L=40.00n
XX0 BA A1 net25 VNW PHVT11LL_CKT W=2.85u L=40.00n
XX2 net25 A2 VDD VNW PHVT11LL_CKT W=2.85u L=40.00n
.ENDS OR4V16_12TH40
.SUBCKT OR4V1RD_12TH40 A1 A2 A3 A4 Z VDD VSS
XX22 DC A4 VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX23 DC A3 VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX19 Z BA net34 VPW NHVT11LL_CKT W=430.00n L=40.00n
XX6 BA A2 VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX5 BA A1 VSS VPW NHVT11LL_CKT W=320.00n L=40.00n
XX18 net34 DC VSS VPW NHVT11LL_CKT W=430.00n L=40.00n
XX20 DC A3 net21 VNW PHVT11LL_CKT W=760.00n L=40.00n
XX21 net21 A4 VDD VNW PHVT11LL_CKT W=760.00n L=40.00n
XX16 Z BA VDD VNW PHVT11LL_CKT W=380.00n L=40.00n
XX17 Z DC VDD VNW PHVT11LL_CKT W=380.00n L=40.00n
XX0 BA A1 net25 VNW PHVT11LL_CKT W=760.00n L=40.00n
XX2 net25 A2 VDD VNW PHVT11LL_CKT W=760.00n L=40.00n
.ENDS OR4V1RD_12TH40
.SUBCKT OR4V1_12TH40 A1 A2 A3 A4 Z VDD VSS
XX22 DC A4 VSS VPW NHVT11LL_CKT W=0.145u L=40.00n
XX23 DC A3 VSS VPW NHVT11LL_CKT W=0.145u L=40.00n
XX19 Z BA net34 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX6 BA A2 VSS VPW NHVT11LL_CKT W=0.145u L=40.00n
XX5 BA A1 VSS VPW NHVT11LL_CKT W=0.145u L=40.00n
XX18 net34 DC VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX20 DC A3 net21 VNW PHVT11LL_CKT W=0.31u L=40.00n
XX21 net21 A4 VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX16 Z BA VDD VNW PHVT11LL_CKT W=0.28u L=40.00n
XX17 Z DC VDD VNW PHVT11LL_CKT W=0.28u L=40.00n
XX0 BA A1 net25 VNW PHVT11LL_CKT W=0.31u L=40.00n
XX2 net25 A2 VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
.ENDS OR4V1_12TH40
.SUBCKT OR4V2RD_12TH40 A1 A2 A3 A4 Z VDD VSS
XX22 DC A4 VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX23 DC A3 VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX19 Z BA net34 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX6 BA A2 VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX5 BA A1 VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX18 net34 DC VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX20 DC A3 net21 VNW PHVT11LL_CKT W=1.08u L=40.00n
XX21 net21 A4 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX16 Z BA VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX17 Z DC VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX0 BA A1 net25 VNW PHVT11LL_CKT W=1.08u L=40.00n
XX2 net25 A2 VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
.ENDS OR4V2RD_12TH40
.SUBCKT OR4V2_12TH40 A1 A2 A3 A4 Z VDD VSS
XX22 DC A4 VSS VPW NHVT11LL_CKT W=185.00n L=40.00n
XX23 DC A3 VSS VPW NHVT11LL_CKT W=185.00n L=40.00n
XX19 Z BA net34 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX6 BA A2 VSS VPW NHVT11LL_CKT W=185.00n L=40.00n
XX5 BA A1 VSS VPW NHVT11LL_CKT W=185.00n L=40.00n
XX18 net34 DC VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX20 DC A3 net21 VNW PHVT11LL_CKT W=395.00n L=40.00n
XX21 net21 A4 VDD VNW PHVT11LL_CKT W=395.00n L=40.00n
XX16 Z BA VDD VNW PHVT11LL_CKT W=395.00n L=40.00n
XX17 Z DC VDD VNW PHVT11LL_CKT W=395.00n L=40.00n
XX0 BA A1 net25 VNW PHVT11LL_CKT W=395.00n L=40.00n
XX2 net25 A2 VDD VNW PHVT11LL_CKT W=395.00n L=40.00n
.ENDS OR4V2_12TH40
.SUBCKT OR4V3_12TH40 A1 A2 A3 A4 Z VDD VSS
XX22 DC A4 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX23 DC A3 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX19 Z BA net34 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX6 BA A2 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX5 BA A1 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX18 net34 DC VSS VPW NHVT11LL_CKT W=0.86u L=40.00n
XX20 DC A3 net21 VNW PHVT11LL_CKT W=0.525u L=40.00n
XX21 net21 A4 VDD VNW PHVT11LL_CKT W=0.525u L=40.00n
XX16 Z BA VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX17 Z DC VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX0 BA A1 net25 VNW PHVT11LL_CKT W=0.525u L=40.00n
XX2 net25 A2 VDD VNW PHVT11LL_CKT W=0.525u L=40.00n
.ENDS OR4V3_12TH40
.SUBCKT OR4V4RD_12TH40 A1 A2 A3 A4 Z VDD VSS
XX22 DC A4 VSS VPW NHVT11LL_CKT W=800.00n L=40.00n
XX23 DC A3 VSS VPW NHVT11LL_CKT W=800.00n L=40.00n
XX19 Z BA net34 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX6 BA A2 VSS VPW NHVT11LL_CKT W=800.00n L=40.00n
XX5 BA A1 VSS VPW NHVT11LL_CKT W=800.00n L=40.00n
XX18 net34 DC VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX20 DC A3 net21 VNW PHVT11LL_CKT W=2.16u L=40.00n
XX21 net21 A4 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
XX16 Z BA VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX17 Z DC VDD VNW PHVT11LL_CKT W=1.08u L=40.00n
XX0 BA A1 net25 VNW PHVT11LL_CKT W=2.16u L=40.00n
XX2 net25 A2 VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
.ENDS OR4V4RD_12TH40
.SUBCKT OR4V4_12TH40 A1 A2 A3 A4 Z VDD VSS
XX22 DC A4 VSS VPW NHVT11LL_CKT W=0.36u L=40.00n
XX23 DC A3 VSS VPW NHVT11LL_CKT W=0.36u L=40.00n
XX19 Z BA net34 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX6 BA A2 VSS VPW NHVT11LL_CKT W=0.36u L=40.00n
XX5 BA A1 VSS VPW NHVT11LL_CKT W=0.36u L=40.00n
XX18 net34 DC VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX20 DC A3 net21 VNW PHVT11LL_CKT W=0.76u L=40.00n
XX21 net21 A4 VDD VNW PHVT11LL_CKT W=0.76u L=40.00n
XX16 Z BA VDD VNW PHVT11LL_CKT W=0.79u L=40.00n
XX17 Z DC VDD VNW PHVT11LL_CKT W=0.79u L=40.00n
XX0 BA A1 net25 VNW PHVT11LL_CKT W=0.76u L=40.00n
XX2 net25 A2 VDD VNW PHVT11LL_CKT W=0.76u L=40.00n
.ENDS OR4V4_12TH40
.SUBCKT OR4V6RD_12TH40 A1 A2 A3 A4 Z VDD VSS
XX22 DC A4 VSS VPW NHVT11LL_CKT W=1.2u L=40.00n
XX23 DC A3 VSS VPW NHVT11LL_CKT W=1.2u L=40.00n
XX19 Z BA net34 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX6 BA A2 VSS VPW NHVT11LL_CKT W=1.2u L=40.00n
XX5 BA A1 VSS VPW NHVT11LL_CKT W=1.2u L=40.00n
XX18 net34 DC VSS VPW NHVT11LL_CKT W=1.83u L=40.00n
XX20 DC A3 net21 VNW PHVT11LL_CKT W=3.24u L=40.00n
XX21 net21 A4 VDD VNW PHVT11LL_CKT W=3.24u L=40.00n
XX16 Z BA VDD VNW PHVT11LL_CKT W=1.62u L=40.00n
XX17 Z DC VDD VNW PHVT11LL_CKT W=1.62u L=40.00n
XX0 BA A1 net25 VNW PHVT11LL_CKT W=3.24u L=40.00n
XX2 net25 A2 VDD VNW PHVT11LL_CKT W=3.24u L=40.00n
.ENDS OR4V6RD_12TH40
.SUBCKT OR4V6_12TH40 A1 A2 A3 A4 Z VDD VSS
XX22 DC A4 VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX23 DC A3 VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX19 Z BA net34 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX6 BA A2 VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX5 BA A1 VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX18 net34 DC VSS VPW NHVT11LL_CKT W=1.83u L=40.00n
XX20 DC A3 net21 VNW PHVT11LL_CKT W=1.07u L=40.00n
XX21 net21 A4 VDD VNW PHVT11LL_CKT W=1.07u L=40.00n
XX16 Z BA VDD VNW PHVT11LL_CKT W=1.185u L=40.00n
XX17 Z DC VDD VNW PHVT11LL_CKT W=1.185u L=40.00n
XX0 BA A1 net25 VNW PHVT11LL_CKT W=1.07u L=40.00n
XX2 net25 A2 VDD VNW PHVT11LL_CKT W=1.07u L=40.00n
.ENDS OR4V6_12TH40
.SUBCKT OR4V8RD_12TH40 A1 A2 A3 A4 Z VDD VSS
XX22 DC A4 VSS VPW NHVT11LL_CKT W=1.6u L=40.00n
XX23 DC A3 VSS VPW NHVT11LL_CKT W=1.6u L=40.00n
XX19 Z BA net34 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX6 BA A2 VSS VPW NHVT11LL_CKT W=1.6u L=40.00n
XX5 BA A1 VSS VPW NHVT11LL_CKT W=1.6u L=40.00n
XX18 net34 DC VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX20 DC A3 net21 VNW PHVT11LL_CKT W=4.34u L=40.00n
XX21 net21 A4 VDD VNW PHVT11LL_CKT W=4.34u L=40.00n
XX16 Z BA VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
XX17 Z DC VDD VNW PHVT11LL_CKT W=2.16u L=40.00n
XX0 BA A1 net25 VNW PHVT11LL_CKT W=4.34u L=40.00n
XX2 net25 A2 VDD VNW PHVT11LL_CKT W=4.34u L=40.00n
.ENDS OR4V8RD_12TH40
.SUBCKT OR4V8_12TH40 A1 A2 A3 A4 Z VDD VSS
XX22 DC A4 VSS VPW NHVT11LL_CKT W=0.69u L=40.00n
XX23 DC A3 VSS VPW NHVT11LL_CKT W=0.69u L=40.00n
XX19 Z BA net34 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX6 BA A2 VSS VPW NHVT11LL_CKT W=0.69u L=40.00n
XX5 BA A1 VSS VPW NHVT11LL_CKT W=0.69u L=40.00n
XX18 net34 DC VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX20 DC A3 net21 VNW PHVT11LL_CKT W=1.455u L=40.00n
XX21 net21 A4 VDD VNW PHVT11LL_CKT W=1.455u L=40.00n
XX16 Z BA VDD VNW PHVT11LL_CKT W=1.58u L=40.00n
XX17 Z DC VDD VNW PHVT11LL_CKT W=1.58u L=40.00n
XX0 BA A1 net25 VNW PHVT11LL_CKT W=1.455u L=40.00n
XX2 net25 A2 VDD VNW PHVT11LL_CKT W=1.455u L=40.00n
.ENDS OR4V8_12TH40
.SUBCKT OR6V0_12TH40 A1 A2 A3 A4 A5 A6 Z VDD VSS
XX4 CBA A3 VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX3 FED A6 VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX5 CBA A1 VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX6 CBA A2 VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX22 FED A5 VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX23 FED A4 VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX18 net31 FED VSS VPW NHVT11LL_CKT W=0.305u L=40.00n
XX19 Z CBA net31 VPW NHVT11LL_CKT W=0.305u L=40.00n
XX7 net58 A3 VDD VNW PHVT11LL_CKT W=0.47u L=40.00n
XX1 net54 A6 VDD VNW PHVT11LL_CKT W=0.47u L=40.00n
XX2 net62 A2 net58 VNW PHVT11LL_CKT W=0.47u L=40.00n
XX0 CBA A1 net62 VNW PHVT11LL_CKT W=0.47u L=40.00n
XX20 FED A4 net50 VNW PHVT11LL_CKT W=0.47u L=40.00n
XX21 net50 A5 net54 VNW PHVT11LL_CKT W=0.47u L=40.00n
XX16 Z CBA VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX17 Z FED VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
.ENDS OR6V0_12TH40
.SUBCKT OR6V12_12TH40 A1 A2 A3 A4 A5 A6 Z VDD VSS
XX4 CBA A3 VSS VPW NHVT11LL_CKT W=1.33u L=40.00n
XX3 FED A6 VSS VPW NHVT11LL_CKT W=1.33u L=40.00n
XX5 CBA A1 VSS VPW NHVT11LL_CKT W=1.33u L=40.00n
XX6 CBA A2 VSS VPW NHVT11LL_CKT W=1.33u L=40.00n
XX22 FED A5 VSS VPW NHVT11LL_CKT W=1.33u L=40.00n
XX23 FED A4 VSS VPW NHVT11LL_CKT W=1.33u L=40.00n
XX18 net31 FED VSS VPW NHVT11LL_CKT W=3.66u L=40.00n
XX19 Z CBA net31 VPW NHVT11LL_CKT W=3.66u L=40.00n
XX7 net58 A3 VDD VNW PHVT11LL_CKT W=4.025u L=40.00n
XX1 net54 A6 VDD VNW PHVT11LL_CKT W=4.025u L=40.00n
XX2 net62 A2 net58 VNW PHVT11LL_CKT W=4.025u L=40.00n
XX0 CBA A1 net62 VNW PHVT11LL_CKT W=4.025u L=40.00n
XX20 FED A4 net50 VNW PHVT11LL_CKT W=4.025u L=40.00n
XX21 net50 A5 net54 VNW PHVT11LL_CKT W=4.025u L=40.00n
XX16 Z CBA VDD VNW PHVT11LL_CKT W=2.37u L=40.00n
XX17 Z FED VDD VNW PHVT11LL_CKT W=2.37u L=40.00n
.ENDS OR6V12_12TH40
.SUBCKT OR6V1_12TH40 A1 A2 A3 A4 A5 A6 Z VDD VSS
XX4 CBA A3 VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX3 FED A6 VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX5 CBA A1 VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX6 CBA A2 VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX22 FED A5 VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX23 FED A4 VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX18 net31 FED VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX19 Z CBA net31 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX7 net58 A3 VDD VNW PHVT11LL_CKT W=0.565u L=40.00n
XX1 net54 A6 VDD VNW PHVT11LL_CKT W=0.565u L=40.00n
XX2 net62 A2 net58 VNW PHVT11LL_CKT W=0.565u L=40.00n
XX0 CBA A1 net62 VNW PHVT11LL_CKT W=0.565u L=40.00n
XX20 FED A4 net50 VNW PHVT11LL_CKT W=0.565u L=40.00n
XX21 net50 A5 net54 VNW PHVT11LL_CKT W=0.565u L=40.00n
XX16 Z CBA VDD VNW PHVT11LL_CKT W=0.28u L=40.00n
XX17 Z FED VDD VNW PHVT11LL_CKT W=0.28u L=40.00n
.ENDS OR6V1_12TH40
.SUBCKT OR6V2_12TH40 A1 A2 A3 A4 A5 A6 Z VDD VSS
XX4 CBA A3 VSS VPW NHVT11LL_CKT W=260.00n L=40.00n
XX3 FED A6 VSS VPW NHVT11LL_CKT W=260.00n L=40.00n
XX5 CBA A1 VSS VPW NHVT11LL_CKT W=260.00n L=40.00n
XX6 CBA A2 VSS VPW NHVT11LL_CKT W=260.00n L=40.00n
XX22 FED A5 VSS VPW NHVT11LL_CKT W=260.00n L=40.00n
XX23 FED A4 VSS VPW NHVT11LL_CKT W=260.00n L=40.00n
XX18 net31 FED VSS VPW NHVT11LL_CKT W=610.00n L=40.00n
XX19 Z CBA net31 VPW NHVT11LL_CKT W=610.00n L=40.00n
XX7 net58 A3 VDD VNW PHVT11LL_CKT W=780.00n L=40.00n
XX1 net54 A6 VDD VNW PHVT11LL_CKT W=780.00n L=40.00n
XX2 net62 A2 net58 VNW PHVT11LL_CKT W=780.00n L=40.00n
XX0 CBA A1 net62 VNW PHVT11LL_CKT W=780.00n L=40.00n
XX20 FED A4 net50 VNW PHVT11LL_CKT W=780.00n L=40.00n
XX21 net50 A5 net54 VNW PHVT11LL_CKT W=780.00n L=40.00n
XX16 Z CBA VDD VNW PHVT11LL_CKT W=395.00n L=40.00n
XX17 Z FED VDD VNW PHVT11LL_CKT W=395.00n L=40.00n
.ENDS OR6V2_12TH40
.SUBCKT OR6V3_12TH40 A1 A2 A3 A4 A5 A6 Z VDD VSS
XX4 CBA A3 VSS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX3 FED A6 VSS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX5 CBA A1 VSS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX6 CBA A2 VSS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX22 FED A5 VSS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX23 FED A4 VSS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX18 net31 FED VSS VPW NHVT11LL_CKT W=0.86u L=40.00n
XX19 Z CBA net31 VPW NHVT11LL_CKT W=0.86u L=40.00n
XX7 net58 A3 VDD VNW PHVT11LL_CKT W=1u L=40.00n
XX1 net54 A6 VDD VNW PHVT11LL_CKT W=1u L=40.00n
XX2 net62 A2 net58 VNW PHVT11LL_CKT W=1u L=40.00n
XX0 CBA A1 net62 VNW PHVT11LL_CKT W=1u L=40.00n
XX20 FED A4 net50 VNW PHVT11LL_CKT W=1u L=40.00n
XX21 net50 A5 net54 VNW PHVT11LL_CKT W=1u L=40.00n
XX16 Z CBA VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX17 Z FED VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
.ENDS OR6V3_12TH40
.SUBCKT OR6V4_12TH40 A1 A2 A3 A4 A5 A6 Z VDD VSS
XX4 CBA A3 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX3 FED A6 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX5 CBA A1 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX6 CBA A2 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX22 FED A5 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX23 FED A4 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX18 net31 FED VSS VPW NHVT11LL_CKT W=1.22u L=40.00n
XX19 Z CBA net31 VPW NHVT11LL_CKT W=1.22u L=40.00n
XX7 net58 A3 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 net54 A6 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX2 net62 A2 net58 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 CBA A1 net62 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX20 FED A4 net50 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX21 net50 A5 net54 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX16 Z CBA VDD VNW PHVT11LL_CKT W=0.79u L=40.00n
XX17 Z FED VDD VNW PHVT11LL_CKT W=0.79u L=40.00n
.ENDS OR6V4_12TH40
.SUBCKT OR6V6_12TH40 A1 A2 A3 A4 A5 A6 Z VDD VSS
XX4 CBA A3 VSS VPW NHVT11LL_CKT W=0.6u L=40.00n
XX3 FED A6 VSS VPW NHVT11LL_CKT W=0.6u L=40.00n
XX5 CBA A1 VSS VPW NHVT11LL_CKT W=0.6u L=40.00n
XX6 CBA A2 VSS VPW NHVT11LL_CKT W=0.6u L=40.00n
XX22 FED A5 VSS VPW NHVT11LL_CKT W=0.6u L=40.00n
XX23 FED A4 VSS VPW NHVT11LL_CKT W=0.6u L=40.00n
XX18 net31 FED VSS VPW NHVT11LL_CKT W=1.83u L=40.00n
XX19 Z CBA net31 VPW NHVT11LL_CKT W=1.83u L=40.00n
XX7 net58 A3 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX1 net54 A6 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX2 net62 A2 net58 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX0 CBA A1 net62 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX20 FED A4 net50 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX21 net50 A5 net54 VNW PHVT11LL_CKT W=1.83u L=40.00n
XX16 Z CBA VDD VNW PHVT11LL_CKT W=1.185u L=40.00n
XX17 Z FED VDD VNW PHVT11LL_CKT W=1.185u L=40.00n
.ENDS OR6V6_12TH40
.SUBCKT OR6V8_12TH40 A1 A2 A3 A4 A5 A6 Z VDD VSS
XX4 CBA A3 VSS VPW NHVT11LL_CKT W=0.8u L=40.00n
XX3 FED A6 VSS VPW NHVT11LL_CKT W=0.8u L=40.00n
XX5 CBA A1 VSS VPW NHVT11LL_CKT W=0.8u L=40.00n
XX6 CBA A2 VSS VPW NHVT11LL_CKT W=0.8u L=40.00n
XX22 FED A5 VSS VPW NHVT11LL_CKT W=0.8u L=40.00n
XX23 FED A4 VSS VPW NHVT11LL_CKT W=0.8u L=40.00n
XX18 net31 FED VSS VPW NHVT11LL_CKT W=2.44u L=40.00n
XX19 Z CBA net31 VPW NHVT11LL_CKT W=2.44u L=40.00n
XX7 net58 A3 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX1 net54 A6 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX2 net62 A2 net58 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX0 CBA A1 net62 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX20 FED A4 net50 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX21 net50 A5 net54 VNW PHVT11LL_CKT W=2.44u L=40.00n
XX16 Z CBA VDD VNW PHVT11LL_CKT W=1.58u L=40.00n
XX17 Z FED VDD VNW PHVT11LL_CKT W=1.58u L=40.00n
.ENDS OR6V8_12TH40
.SUBCKT PULL0_12TH40 Z VDD VSS
XX0 Z net4 VSS VPW NHVT11LL_CKT W=560.00n L=40.00n
XX2 net2 net4 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX1 net4 net2 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX3 net4 net4 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS PULL0_12TH40
.SUBCKT PULL1_12TH40 Z VDD VSS
XX2 net8 net6 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX0 net8 net8 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX1 net6 net8 VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX3 Z net8 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS PULL1_12TH40
.SUBCKT SDGRNQNV2_12TH40 CK D QN RN SE SI VDD VSS
XX0 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX5 net83 D net15 VPW NHVT11LL_CKT W=0.405u L=40.00n
XX6 net15 RN net19 VPW NHVT11LL_CKT W=0.5u L=40.00n
XX7 net19 SEN VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX10 net23 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX11 net83 SE net23 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX13 net83 cn net34 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX15 net35 net34 VSS VPW NHVT11LL_CKT W=0.475u L=40.00n
XX17 net39 net35 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX19 net34 c net39 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX21 net35 c net50 VPW NHVT11LL_CKT W=0.39u L=40.00n
XX27 net51 net50 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net50 cn net59 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net59 net51 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 QN net50 VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX31 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX1 SEN SE VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX2 net86 SE VDD VNW PHVT11LL_CKT W=0.555u L=40.00n
XX3 net83 D net86 VNW PHVT11LL_CKT W=0.405u L=40.00n
XX4 net83 RN net86 VNW PHVT11LL_CKT W=0.25u L=40.00n
XX9 net98 SI VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX8 net83 SEN net98 VNW PHVT11LL_CKT W=0.14u L=40.00n
XX12 net83 c net34 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX14 net35 net34 VDD VNW PHVT11LL_CKT W=0.495u L=40.00n
XX16 net114 net35 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX18 net34 cn net114 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 net126 net51 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 net51 net50 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX22 net50 c net126 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net35 cn net50 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX28 QN net50 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX32 c cn VDD VNW PHVT11LL_CKT W=0.45u L=40.00n
XX30 cn CK VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS SDGRNQNV2_12TH40
.SUBCKT SDGRNQNV4_12TH40 CK D QN RN SE SI VDD VSS
XX0 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX5 net83 D net15 VPW NHVT11LL_CKT W=0.405u L=40.00n
XX6 net15 RN net19 VPW NHVT11LL_CKT W=0.5u L=40.00n
XX7 net19 SEN VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX10 net23 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX11 net83 SE net23 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX13 net83 cn net34 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX15 net35 net34 VSS VPW NHVT11LL_CKT W=0.475u L=40.00n
XX17 net39 net35 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX19 net34 c net39 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX21 net35 c net50 VPW NHVT11LL_CKT W=0.39u L=40.00n
XX27 net51 net50 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net50 cn net59 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net59 net51 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 QN net50 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX31 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX33 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX1 SEN SE VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX2 net86 SE VDD VNW PHVT11LL_CKT W=0.555u L=40.00n
XX3 net83 D net86 VNW PHVT11LL_CKT W=0.465u L=40.00n
XX4 net83 RN net86 VNW PHVT11LL_CKT W=0.25u L=40.00n
XX9 net98 SI VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX8 net83 SEN net98 VNW PHVT11LL_CKT W=0.14u L=40.00n
XX12 net83 c net34 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX14 net35 net34 VDD VNW PHVT11LL_CKT W=0.565u L=40.00n
XX16 net114 net35 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX18 net34 cn net114 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 net126 net51 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 net51 net50 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX22 net50 c net126 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net35 cn net50 VNW PHVT11LL_CKT W=0.4u L=40.00n
XX28 QN net50 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX32 c cn VDD VNW PHVT11LL_CKT W=0.38u L=40.00n
XX30 cn CK VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
.ENDS SDGRNQNV4_12TH40
.SUBCKT SDGRNQNV6_12TH40 CK D QN RN SE SI VDD VSS
XX0 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX5 net83 D net15 VPW NHVT11LL_CKT W=0.42u L=40.00n
XX6 net15 RN net19 VPW NHVT11LL_CKT W=0.5u L=40.00n
XX7 net19 SEN VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX10 net23 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX11 net83 SE net23 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX13 net83 cn net34 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX15 net35 net34 VSS VPW NHVT11LL_CKT W=0.56u L=40.00n
XX17 net39 net35 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX19 net34 c net39 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX21 net35 c net50 VPW NHVT11LL_CKT W=0.44u L=40.00n
XX27 net51 net50 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net50 cn net59 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net59 net51 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 QN net50 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX31 cn CK VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX33 c cn VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX1 SEN SE VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX2 net86 SE VDD VNW PHVT11LL_CKT W=0.57u L=40.00n
XX3 net83 D net86 VNW PHVT11LL_CKT W=0.57u L=40.00n
XX4 net83 RN net86 VNW PHVT11LL_CKT W=0.25u L=40.00n
XX9 net98 SI VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX8 net83 SEN net98 VNW PHVT11LL_CKT W=0.14u L=40.00n
XX12 net83 c net34 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX14 net35 net34 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX16 net114 net35 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX18 net34 cn net114 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 net126 net51 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 net51 net50 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX22 net50 c net126 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net35 cn net50 VNW PHVT11LL_CKT W=0.49u L=40.00n
XX28 QN net50 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX32 c cn VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX30 cn CK VDD VNW PHVT11LL_CKT W=0.21u L=40.00n
.ENDS SDGRNQNV6_12TH40
.SUBCKT SDGRNQV2_12TH40 CK D Q RN SE SI VDD VSS
XX0 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX5 net83 D net15 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX6 net15 RN net19 VPW NHVT11LL_CKT W=0.5u L=40.00n
XX7 net19 SEN VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX10 net23 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX11 net83 SE net23 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX13 net83 cn net34 VPW NHVT11LL_CKT W=0.26u L=40.00n
XX15 net35 net34 VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX17 net39 net35 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX19 net34 c net39 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX21 net35 c net50 VPW NHVT11LL_CKT W=0.26u L=40.00n
XX27 net51 net50 VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX26 net50 cn net59 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net59 net51 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 Q net51 VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX31 cn CK VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX33 c cn VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX1 SEN SE VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX2 net86 SE VDD VNW PHVT11LL_CKT W=0.58u L=40.00n
XX3 net83 D net86 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX4 net83 RN net86 VNW PHVT11LL_CKT W=0.25u L=40.00n
XX9 net98 SI VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX8 net83 SEN net98 VNW PHVT11LL_CKT W=0.14u L=40.00n
XX12 net83 c net34 VNW PHVT11LL_CKT W=0.26u L=40.00n
XX14 net35 net34 VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX16 net114 net35 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX18 net34 cn net114 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 net126 net51 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 net51 net50 VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX22 net50 c net126 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net35 cn net50 VNW PHVT11LL_CKT W=0.28u L=40.00n
XX28 Q net51 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX32 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX30 cn CK VDD VNW PHVT11LL_CKT W=0.13u L=40.00n
.ENDS SDGRNQV2_12TH40
.SUBCKT SDGRNQV4_12TH40 CK D Q RN SE SI VDD VSS
XX0 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX5 net83 D net15 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX6 net15 RN net19 VPW NHVT11LL_CKT W=0.5u L=40.00n
XX7 net19 SEN VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX10 net23 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX11 net83 SE net23 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX13 net83 cn net34 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX15 net35 net34 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX17 net39 net35 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX19 net34 c net39 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX21 net35 c net50 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX27 net51 net50 VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX26 net50 cn net59 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net59 net51 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 Q net51 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX31 cn CK VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX33 c cn VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX1 SEN SE VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX2 net86 SE VDD VNW PHVT11LL_CKT W=0.58u L=40.00n
XX3 net83 D net86 VNW PHVT11LL_CKT W=0.49u L=40.00n
XX4 net83 RN net86 VNW PHVT11LL_CKT W=0.25u L=40.00n
XX9 net98 SI VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX8 net83 SEN net98 VNW PHVT11LL_CKT W=0.14u L=40.00n
XX12 net83 c net34 VNW PHVT11LL_CKT W=0.34u L=40.00n
XX14 net35 net34 VDD VNW PHVT11LL_CKT W=0.48u L=40.00n
XX16 net114 net35 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX18 net34 cn net114 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 net126 net51 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 net51 net50 VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX22 net50 c net126 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net35 cn net50 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX28 Q net51 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX32 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX30 cn CK VDD VNW PHVT11LL_CKT W=0.18u L=40.00n
.ENDS SDGRNQV4_12TH40
.SUBCKT SDGRNQV6_12TH40 CK D Q RN SE SI VDD VSS
XX0 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX5 net83 D net15 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX6 net15 RN net19 VPW NHVT11LL_CKT W=0.5u L=40.00n
XX7 net19 SEN VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX10 net23 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX11 net83 SE net23 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX13 net83 cn net34 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX15 net35 net34 VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX17 net39 net35 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX19 net34 c net39 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX21 net35 c net50 VPW NHVT11LL_CKT W=0.42u L=40.00n
XX27 net51 net50 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX26 net50 cn net59 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net59 net51 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 Q net51 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX31 cn CK VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX33 c cn VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX1 SEN SE VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX2 net86 SE VDD VNW PHVT11LL_CKT W=0.58u L=40.00n
XX3 net83 D net86 VNW PHVT11LL_CKT W=0.58u L=40.00n
XX4 net83 RN net86 VNW PHVT11LL_CKT W=0.25u L=40.00n
XX9 net98 SI VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX8 net83 SEN net98 VNW PHVT11LL_CKT W=0.14u L=40.00n
XX12 net83 c net34 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX14 net35 net34 VDD VNW PHVT11LL_CKT W=0.49u L=40.00n
XX16 net114 net35 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX18 net34 cn net114 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 net126 net51 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 net51 net50 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX22 net50 c net126 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net35 cn net50 VNW PHVT11LL_CKT W=0.35u L=40.00n
XX28 Q net51 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX32 c cn VDD VNW PHVT11LL_CKT W=0.47u L=40.00n
XX30 cn CK VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
.ENDS SDGRNQV6_12TH40
.SUBCKT SDGRSNQNV2_12TH40 CK D QN RN SE SI SN VDD VSS
XX17 net140 cn M VPW NHVT11LL_CKT W=0.33u L=40.00n
XX29 S c OS VPW NHVT11LL_CKT W=0.37u L=40.00n
XX37 VSS net112 net95 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX36 net95 cn OS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 VSS S net103 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX24 net103 c M VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 QN OS VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX31 net112 OS VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX21 S M VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX27 SEN SE VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX19 SNN SN VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX15 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX11 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net136 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX8 net140 SE net136 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX5 net144 SEN VSS VPW NHVT11LL_CKT W=0.48u L=40.00n
XX13 net140 SNN net152 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX4 net152 RN net144 VPW NHVT11LL_CKT W=0.48u L=40.00n
XX3 net140 D net152 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX16 net140 c M VNW PHVT11LL_CKT W=0.495u L=40.00n
XX28 S cn OS VNW PHVT11LL_CKT W=0.33u L=40.00n
XX35 net16 c OS VNW PHVT11LL_CKT W=120.00n L=40.00n
XX34 VDD net112 net16 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 net24 cn M VNW PHVT11LL_CKT W=120.00n L=40.00n
XX22 VDD S net24 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX32 QN OS VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX30 net112 OS VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX26 SEN SE VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX18 SNN SN VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX14 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX10 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX20 S M VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX7 net140 SEN net63 VNW PHVT11LL_CKT W=0.14u L=40.00n
XX6 net63 SI VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX2 net140 D net71 VNW PHVT11LL_CKT W=0.6u L=40.00n
XX1 net71 SNN net75 VNW PHVT11LL_CKT W=0.6u L=40.00n
XX12 net140 RN net75 VNW PHVT11LL_CKT W=0.25u L=40.00n
XX0 net75 SE VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
.ENDS SDGRSNQNV2_12TH40
.SUBCKT SDGRSNQNV4_12TH40 CK D QN RN SE SI SN VDD VSS
XX17 net140 cn M VPW NHVT11LL_CKT W=0.33u L=40.00n
XX29 S c OS VPW NHVT11LL_CKT W=0.37u L=40.00n
XX37 VSS net112 net95 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX36 net95 cn OS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 VSS S net103 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX24 net103 c M VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 QN OS VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX31 net112 OS VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX21 S M VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX27 SEN SE VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX19 SNN SN VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX15 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX11 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net136 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX8 net140 SE net136 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX5 net144 SEN VSS VPW NHVT11LL_CKT W=0.48u L=40.00n
XX13 net140 SNN net152 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX4 net152 RN net144 VPW NHVT11LL_CKT W=0.48u L=40.00n
XX3 net140 D net152 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX16 net140 c M VNW PHVT11LL_CKT W=0.495u L=40.00n
XX28 S cn OS VNW PHVT11LL_CKT W=0.37u L=40.00n
XX35 net16 c OS VNW PHVT11LL_CKT W=120.00n L=40.00n
XX34 VDD net112 net16 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 net24 cn M VNW PHVT11LL_CKT W=120.00n L=40.00n
XX22 VDD S net24 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX32 QN OS VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX30 net112 OS VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX26 SEN SE VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX18 SNN SN VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX14 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX10 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX20 S M VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX7 net140 SEN net63 VNW PHVT11LL_CKT W=0.14u L=40.00n
XX6 net63 SI VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX2 net140 D net71 VNW PHVT11LL_CKT W=0.6u L=40.00n
XX1 net71 SNN net75 VNW PHVT11LL_CKT W=0.6u L=40.00n
XX12 net140 RN net75 VNW PHVT11LL_CKT W=0.25u L=40.00n
XX0 net75 SE VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
.ENDS SDGRSNQNV4_12TH40
.SUBCKT SDGRSNQNV6_12TH40 CK D QN RN SE SI SN VDD VSS
XX17 net140 cn M VPW NHVT11LL_CKT W=0.33u L=40.00n
XX29 S c OS VPW NHVT11LL_CKT W=0.37u L=40.00n
XX37 VSS net112 net95 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX36 net95 cn OS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 VSS S net103 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX24 net103 c M VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 QN OS VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX31 net112 OS VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX21 S M VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX27 SEN SE VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX19 SNN SN VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX15 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX11 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net136 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX8 net140 SE net136 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX5 net144 SEN VSS VPW NHVT11LL_CKT W=0.48u L=40.00n
XX13 net140 SNN net152 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX4 net152 RN net144 VPW NHVT11LL_CKT W=0.48u L=40.00n
XX3 net140 D net152 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX16 net140 c M VNW PHVT11LL_CKT W=0.495u L=40.00n
XX28 S cn OS VNW PHVT11LL_CKT W=0.45u L=40.00n
XX35 net16 c OS VNW PHVT11LL_CKT W=120.00n L=40.00n
XX34 VDD net112 net16 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 net24 cn M VNW PHVT11LL_CKT W=120.00n L=40.00n
XX22 VDD S net24 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX32 QN OS VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX30 net112 OS VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX26 SEN SE VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX18 SNN SN VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX14 c cn VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX10 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX20 S M VDD VNW PHVT11LL_CKT W=0.605u L=40.00n
XX7 net140 SEN net63 VNW PHVT11LL_CKT W=0.14u L=40.00n
XX6 net63 SI VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX2 net140 D net71 VNW PHVT11LL_CKT W=0.6u L=40.00n
XX1 net71 SNN net75 VNW PHVT11LL_CKT W=0.6u L=40.00n
XX12 net140 RN net75 VNW PHVT11LL_CKT W=0.25u L=40.00n
XX0 net75 SE VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
.ENDS SDGRSNQNV6_12TH40
.SUBCKT SDGRSNQV2_12TH40 CK D Q RN SE SI SN VDD VSS
XX17 net140 cn M VPW NHVT11LL_CKT W=0.33u L=40.00n
XX29 S c OS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX37 VSS net112 net95 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX36 net95 cn OS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 VSS S net103 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX24 net103 c M VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 Q net112 VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX31 net112 OS VSS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX21 S M VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX27 SEN SE VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX19 SNN SN VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX15 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX11 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net136 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX8 net140 SE net136 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX5 net144 SEN VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX13 net140 SNN net152 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX4 net152 RN net144 VPW NHVT11LL_CKT W=0.47u L=40.00n
XX3 net140 D net152 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX16 net140 c M VNW PHVT11LL_CKT W=0.375u L=40.00n
XX28 S cn OS VNW PHVT11LL_CKT W=0.33u L=40.00n
XX35 net16 c OS VNW PHVT11LL_CKT W=120.00n L=40.00n
XX34 VDD net112 net16 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 net24 cn M VNW PHVT11LL_CKT W=120.00n L=40.00n
XX22 VDD S net24 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX32 Q net112 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX30 net112 OS VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX26 SEN SE VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX18 SNN SN VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX14 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX10 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX20 S M VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX7 net140 SEN net63 VNW PHVT11LL_CKT W=0.14u L=40.00n
XX6 net63 SI VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX2 net140 D net71 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX1 net71 SNN net75 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX12 net140 RN net75 VNW PHVT11LL_CKT W=0.25u L=40.00n
XX0 net75 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
.ENDS SDGRSNQV2_12TH40
.SUBCKT SDGRSNQV4_12TH40 CK D Q RN SE SI SN VDD VSS
XX17 net140 cn M VPW NHVT11LL_CKT W=0.33u L=40.00n
XX29 S c OS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX37 VSS net112 net95 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX36 net95 cn OS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 VSS S net103 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX24 net103 c M VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 Q net112 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX31 net112 OS VSS VPW NHVT11LL_CKT W=0.36u L=40.00n
XX21 S M VSS VPW NHVT11LL_CKT W=0.495u L=40.00n
XX27 SEN SE VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX19 SNN SN VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX15 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX11 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net136 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX8 net140 SE net136 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX5 net144 SEN VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX13 net140 SNN net152 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX4 net152 RN net144 VPW NHVT11LL_CKT W=0.47u L=40.00n
XX3 net140 D net152 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX16 net140 c M VNW PHVT11LL_CKT W=0.375u L=40.00n
XX28 S cn OS VNW PHVT11LL_CKT W=0.33u L=40.00n
XX35 net16 c OS VNW PHVT11LL_CKT W=120.00n L=40.00n
XX34 VDD net112 net16 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 net24 cn M VNW PHVT11LL_CKT W=120.00n L=40.00n
XX22 VDD S net24 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX32 Q net112 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX30 net112 OS VDD VNW PHVT11LL_CKT W=0.51u L=40.00n
XX26 SEN SE VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX18 SNN SN VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX14 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX10 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX20 S M VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX7 net140 SEN net63 VNW PHVT11LL_CKT W=0.14u L=40.00n
XX6 net63 SI VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX2 net140 D net71 VNW PHVT11LL_CKT W=0.535u L=40.00n
XX1 net71 SNN net75 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX12 net140 RN net75 VNW PHVT11LL_CKT W=0.25u L=40.00n
XX0 net75 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
.ENDS SDGRSNQV4_12TH40
.SUBCKT SDGRSNQV6_12TH40 CK D Q RN SE SI SN VDD VSS
XX17 net140 cn M VPW NHVT11LL_CKT W=0.33u L=40.00n
XX29 S c OS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX37 VSS net112 net95 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX36 net95 cn OS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 VSS S net103 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX24 net103 c M VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 Q net112 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX31 net112 OS VSS VPW NHVT11LL_CKT W=0.41u L=40.00n
XX21 S M VSS VPW NHVT11LL_CKT W=0.495u L=40.00n
XX27 SEN SE VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX19 SNN SN VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX15 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX11 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net136 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX8 net140 SE net136 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX5 net144 SEN VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX13 net140 SNN net152 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX4 net152 RN net144 VPW NHVT11LL_CKT W=0.47u L=40.00n
XX3 net140 D net152 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX16 net140 c M VNW PHVT11LL_CKT W=0.375u L=40.00n
XX28 S cn OS VNW PHVT11LL_CKT W=0.33u L=40.00n
XX35 net16 c OS VNW PHVT11LL_CKT W=120.00n L=40.00n
XX34 VDD net112 net16 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 net24 cn M VNW PHVT11LL_CKT W=120.00n L=40.00n
XX22 VDD S net24 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX32 Q net112 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX30 net112 OS VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX26 SEN SE VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX18 SNN SN VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX14 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX10 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX20 S M VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX7 net140 SEN net63 VNW PHVT11LL_CKT W=0.14u L=40.00n
XX6 net63 SI VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX2 net140 D net71 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX1 net71 SNN net75 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX12 net140 RN net75 VNW PHVT11LL_CKT W=0.25u L=40.00n
XX0 net75 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
.ENDS SDGRSNQV6_12TH40
.SUBCKT SDGSNQNV2_12TH40 CK D QN SE SI SN VDD VSS
XX12 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX8 net83 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX36 VSS net107 net90 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX35 net90 cn PS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX21 net146 c PM VPW NHVT11LL_CKT W=120.00n L=40.00n
XX32 QN PS VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX26 M c PS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX30 net107 PS VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 M PM VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX16 N74 cn PM VPW NHVT11LL_CKT W=0.33u L=40.00n
XX3 N74 D net123 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX4 net123 SEN VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX24 SNN SN VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX28 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 N74 SE net83 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 N74 SNN net123 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX22 VSS M net146 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX20 net7 cn PM VNW PHVT11LL_CKT W=120.00n L=40.00n
XX34 net11 c PS VNW PHVT11LL_CKT W=120.00n L=40.00n
XX33 VDD net107 net11 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX31 QN PS VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX19 VDD M net7 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX29 net107 PS VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 N74 c PM VNW PHVT11LL_CKT W=330.00n L=40.00n
XX17 M PM VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX2 N74 D net42 VNW PHVT11LL_CKT W=0.44u L=40.00n
XX1 net42 SNN net46 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net46 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX6 N74 SEN net54 VNW PHVT11LL_CKT W=0.14u L=40.00n
XX5 net54 SI VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX27 SEN SE VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX23 SNN SN VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX25 M cn PS VNW PHVT11LL_CKT W=0.33u L=40.00n
.ENDS SDGSNQNV2_12TH40
.SUBCKT SDGSNQNV4_12TH40 CK D QN SE SI SN VDD VSS
XX12 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX8 net83 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX36 VSS net107 net90 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX35 net90 cn PS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX21 net146 c PM VPW NHVT11LL_CKT W=120.00n L=40.00n
XX32 QN PS VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX26 M c PS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX30 net107 PS VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 M PM VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX16 N74 cn PM VPW NHVT11LL_CKT W=0.33u L=40.00n
XX3 N74 D net123 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX4 net123 SEN VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX24 SNN SN VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX28 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 N74 SE net83 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 N74 SNN net123 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX22 VSS M net146 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX20 net7 cn PM VNW PHVT11LL_CKT W=120.00n L=40.00n
XX34 net11 c PS VNW PHVT11LL_CKT W=120.00n L=40.00n
XX33 VDD net107 net11 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX31 QN PS VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX19 VDD M net7 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX29 net107 PS VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 N74 c PM VNW PHVT11LL_CKT W=330.00n L=40.00n
XX17 M PM VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX2 N74 D net42 VNW PHVT11LL_CKT W=0.53u L=40.00n
XX1 net42 SNN net46 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net46 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX6 N74 SEN net54 VNW PHVT11LL_CKT W=0.14u L=40.00n
XX5 net54 SI VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX27 SEN SE VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX23 SNN SN VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX25 M cn PS VNW PHVT11LL_CKT W=0.425u L=40.00n
.ENDS SDGSNQNV4_12TH40
.SUBCKT SDGSNQNV6_12TH40 CK D QN SE SI SN VDD VSS
XX12 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX8 net83 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX36 VSS net107 net90 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX35 net90 cn PS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX21 net146 c PM VPW NHVT11LL_CKT W=120.00n L=40.00n
XX32 QN PS VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX26 M c PS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX30 net107 PS VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 M PM VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX16 N74 cn PM VPW NHVT11LL_CKT W=0.33u L=40.00n
XX3 N74 D net123 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX4 net123 SEN VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX24 SNN SN VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX28 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 N74 SE net83 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 N74 SNN net123 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX22 VSS M net146 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX20 net7 cn PM VNW PHVT11LL_CKT W=120.00n L=40.00n
XX34 net11 c PS VNW PHVT11LL_CKT W=120.00n L=40.00n
XX33 VDD net107 net11 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX31 QN PS VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX19 VDD M net7 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX29 net107 PS VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 N74 c PM VNW PHVT11LL_CKT W=330.00n L=40.00n
XX17 M PM VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX2 N74 D net42 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX1 net42 SNN net46 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net46 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX6 N74 SEN net54 VNW PHVT11LL_CKT W=0.14u L=40.00n
XX5 net54 SI VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX27 SEN SE VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX23 SNN SN VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX25 M cn PS VNW PHVT11LL_CKT W=0.435u L=40.00n
.ENDS SDGSNQNV6_12TH40
.SUBCKT SDGSNQV2_12TH40 CK D Q SE SI SN VDD VSS
XX12 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX8 net83 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX36 VSS net107 net90 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX35 net90 cn PS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX21 net146 c PM VPW NHVT11LL_CKT W=120.00n L=40.00n
XX32 Q net107 VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX26 M c PS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX30 net107 PS VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX18 M PM VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX16 N74 cn PM VPW NHVT11LL_CKT W=0.33u L=40.00n
XX3 N74 D net123 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX4 net123 SEN VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX24 SNN SN VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX28 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 N74 SE net83 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 N74 SNN net123 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX22 VSS M net146 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX20 net7 cn PM VNW PHVT11LL_CKT W=120.00n L=40.00n
XX34 net11 c PS VNW PHVT11LL_CKT W=120.00n L=40.00n
XX33 VDD net107 net11 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX31 Q net107 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX19 VDD M net7 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX29 net107 PS VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX15 N74 c PM VNW PHVT11LL_CKT W=330.00n L=40.00n
XX17 M PM VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX2 N74 D net42 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX1 net42 SNN net46 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net46 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX6 N74 SEN net54 VNW PHVT11LL_CKT W=0.14u L=40.00n
XX5 net54 SI VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX27 SEN SE VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX23 SNN SN VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX25 M cn PS VNW PHVT11LL_CKT W=0.33u L=40.00n
.ENDS SDGSNQV2_12TH40
.SUBCKT SDGSNQV4_12TH40 CK D Q SE SI SN VDD VSS
XX12 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX8 net83 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX36 VSS net107 net90 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX35 net90 cn PS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX21 net146 c PM VPW NHVT11LL_CKT W=120.00n L=40.00n
XX32 Q net107 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX26 M c PS VPW NHVT11LL_CKT W=0.37u L=40.00n
XX30 net107 PS VSS VPW NHVT11LL_CKT W=0.36u L=40.00n
XX18 M PM VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX16 N74 cn PM VPW NHVT11LL_CKT W=0.33u L=40.00n
XX3 N74 D net123 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX4 net123 SEN VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX24 SNN SN VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX28 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 N74 SE net83 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 N74 SNN net123 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX22 VSS M net146 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX20 net7 cn PM VNW PHVT11LL_CKT W=120.00n L=40.00n
XX34 net11 c PS VNW PHVT11LL_CKT W=120.00n L=40.00n
XX33 VDD net107 net11 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX31 Q net107 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX19 VDD M net7 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX29 net107 PS VDD VNW PHVT11LL_CKT W=0.51u L=40.00n
XX15 N74 c PM VNW PHVT11LL_CKT W=330.00n L=40.00n
XX17 M PM VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX2 N74 D net42 VNW PHVT11LL_CKT W=0.52u L=40.00n
XX1 net42 SNN net46 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net46 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX6 N74 SEN net54 VNW PHVT11LL_CKT W=0.14u L=40.00n
XX5 net54 SI VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX27 SEN SE VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX23 SNN SN VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX25 M cn PS VNW PHVT11LL_CKT W=0.35u L=40.00n
.ENDS SDGSNQV4_12TH40
.SUBCKT SDGSNQV6_12TH40 CK D Q SE SI SN VDD VSS
XX12 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX8 net83 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX36 VSS net107 net90 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX35 net90 cn PS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX21 net146 c PM VPW NHVT11LL_CKT W=120.00n L=40.00n
XX32 Q net107 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX26 M c PS VPW NHVT11LL_CKT W=0.39u L=40.00n
XX30 net107 PS VSS VPW NHVT11LL_CKT W=0.39u L=40.00n
XX18 M PM VSS VPW NHVT11LL_CKT W=0.475u L=40.00n
XX16 N74 cn PM VPW NHVT11LL_CKT W=0.33u L=40.00n
XX3 N74 D net123 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX4 net123 SEN VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX24 SNN SN VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX28 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 N74 SE net83 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 N74 SNN net123 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX22 VSS M net146 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX20 net7 cn PM VNW PHVT11LL_CKT W=120.00n L=40.00n
XX34 net11 c PS VNW PHVT11LL_CKT W=120.00n L=40.00n
XX33 VDD net107 net11 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX31 Q net107 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX19 VDD M net7 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX29 net107 PS VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX15 N74 c PM VNW PHVT11LL_CKT W=330.00n L=40.00n
XX17 M PM VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX2 N74 D net42 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX1 net42 SNN net46 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net46 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX6 N74 SEN net54 VNW PHVT11LL_CKT W=0.14u L=40.00n
XX5 net54 SI VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX27 SEN SE VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX23 SNN SN VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX25 M cn PS VNW PHVT11LL_CKT W=0.35u L=40.00n
.ENDS SDGSNQV6_12TH40
.SUBCKT SDQNV0_12TH40 CK D QN SE SI VDD VSS
XX22 QN net37 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX18 net22 net37 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net37 cn net30 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net30 net22 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net46 c net37 VPW NHVT11LL_CKT W=0.32u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net38 net46 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net53 c net38 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net46 net53 VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX3 net54 cn net53 VPW NHVT11LL_CKT W=0.21u L=40.00n
XX2 net54 D net58 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX25 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net58 SEN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX30 net62 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net54 SE net62 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net37 VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX21 net22 net37 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net37 c net93 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net93 net22 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net46 cn net37 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net109 net46 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net53 cn net109 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net46 net53 VDD VNW PHVT11LL_CKT W=0.39u L=40.00n
XX0 net54 c net53 VNW PHVT11LL_CKT W=0.22u L=40.00n
XX1 net54 D net121 VNW PHVT11LL_CKT W=0.31u L=40.00n
XX29 net54 SEN net125 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX28 net125 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX24 SEN SE VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX27 net121 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
.ENDS SDQNV0_12TH40
.SUBCKT SDQNV2_12TH40 CK D QN SE SI VDD VSS
XX22 QN net37 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX18 net22 net37 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net37 cn net30 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net30 net22 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net46 c net37 VPW NHVT11LL_CKT W=330.00n L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=190.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net38 net46 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net53 c net38 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net46 net53 VSS VPW NHVT11LL_CKT W=455.00n L=40.00n
XX3 net54 cn net53 VPW NHVT11LL_CKT W=330.00n L=40.00n
XX2 net54 D net58 VPW NHVT11LL_CKT W=0.34u L=40.00n
XX25 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net58 SEN VSS VPW NHVT11LL_CKT W=0.6u L=40.00n
XX30 net62 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net54 SE net62 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net37 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX21 net22 net37 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net37 c net93 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net93 net22 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net46 cn net37 VNW PHVT11LL_CKT W=0.31u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net109 net46 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net53 cn net109 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net46 net53 VDD VNW PHVT11LL_CKT W=0.41u L=40.00n
XX0 net54 c net53 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX1 net54 D net121 VNW PHVT11LL_CKT W=0.4u L=40.00n
XX29 net54 SEN net125 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX28 net125 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX24 SEN SE VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX27 net121 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
.ENDS SDQNV2_12TH40
.SUBCKT SDQNV4_12TH40 CK D QN SE SI VDD VSS
XX22 QN net37 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX18 net22 net37 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net37 cn net30 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net30 net22 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net46 c net37 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.155u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX9 net38 net46 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net53 c net38 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net46 net53 VSS VPW NHVT11LL_CKT W=0.46u L=40.00n
XX3 net54 cn net53 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX2 net54 D net58 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX25 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net58 SEN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX30 net62 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net54 SE net62 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net37 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX21 net22 net37 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net37 c net93 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net93 net22 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net46 cn net37 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX8 net109 net46 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net53 cn net109 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net46 net53 VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX0 net54 c net53 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX1 net54 D net121 VNW PHVT11LL_CKT W=0.53u L=40.00n
XX29 net54 SEN net125 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX28 net125 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX24 SEN SE VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX27 net121 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
.ENDS SDQNV4_12TH40
.SUBCKT SDQNV6_12TH40 CK D QN SE SI VDD VSS
XX22 QN net37 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX18 net22 net37 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net37 cn net30 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net30 net22 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net46 c net37 VPW NHVT11LL_CKT W=0.42u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX9 net38 net46 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net53 c net38 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net46 net53 VSS VPW NHVT11LL_CKT W=0.47u L=40.00n
XX3 net54 cn net53 VPW NHVT11LL_CKT W=0.32u L=40.00n
XX2 net54 D net58 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX25 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net58 SEN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX30 net62 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net54 SE net62 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net37 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX21 net22 net37 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net37 c net93 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net93 net22 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net46 cn net37 VNW PHVT11LL_CKT W=0.54u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.21u L=40.00n
XX8 net109 net46 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net53 cn net109 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net46 net53 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net54 c net53 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX1 net54 D net121 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX29 net54 SEN net125 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX28 net125 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX24 SEN SE VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX27 net121 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
.ENDS SDQNV6_12TH40
.SUBCKT SDQV0_12TH40 CK D Q SE SI VDD VSS
XX31 net86 SE net78 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net78 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net82 SEN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX2 net86 D net82 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX3 net86 cn net93 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX4 net94 net93 VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX6 net93 c net102 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net102 net94 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net94 c net109 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX16 net110 net118 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net109 cn net110 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net118 net109 VSS VPW NHVT11LL_CKT W=0.135u L=40.00n
XX25 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX22 Q net118 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX27 net25 SE VDD VNW PHVT11LL_CKT W=0.59u L=40.00n
XX28 net21 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX29 net86 SEN net21 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net86 D net25 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX0 net86 c net93 VNW PHVT11LL_CKT W=0.22u L=40.00n
XX5 net94 net93 VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX7 net93 cn net37 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net37 net94 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net94 cn net109 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX19 net53 net118 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net109 c net53 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX21 net118 net109 VDD VNW PHVT11LL_CKT W=0.24u L=40.00n
XX24 SEN SE VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.38u L=40.00n
XX23 Q net118 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
.ENDS SDQV0_12TH40
.SUBCKT SDQV2_12TH40 CK D Q SE SI VDD VSS
XX31 net86 SE net78 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net78 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net82 SEN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX2 net86 D net82 VPW NHVT11LL_CKT W=0.32u L=40.00n
XX3 net86 cn net93 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX4 net94 net93 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX6 net93 c net102 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net102 net94 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net94 c net109 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX16 net110 net118 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net109 cn net110 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net118 net109 VSS VPW NHVT11LL_CKT W=230.00n L=40.00n
XX25 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=130.00n L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=185.00n L=40.00n
XX22 Q net118 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX27 net25 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX28 net21 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX29 net86 SEN net21 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net86 D net25 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX0 net86 c net93 VNW PHVT11LL_CKT W=260.00n L=40.00n
XX5 net94 net93 VDD VNW PHVT11LL_CKT W=440.00n L=40.00n
XX7 net93 cn net37 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net37 net94 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net94 cn net109 VNW PHVT11LL_CKT W=260.00n L=40.00n
XX19 net53 net118 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net109 c net53 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX21 net118 net109 VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX24 SEN SE VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX23 Q net118 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS SDQV2_12TH40
.SUBCKT SDQV4_12TH40 CK D Q SE SI VDD VSS
XX31 net86 SE net78 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net78 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net82 SEN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX2 net86 D net82 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX3 net86 cn net93 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX4 net94 net93 VSS VPW NHVT11LL_CKT W=0.445u L=40.00n
XX6 net93 c net102 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net102 net94 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net94 c net109 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX16 net110 net118 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net109 cn net110 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net118 net109 VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX25 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX22 Q net118 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX27 net25 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX28 net21 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX29 net86 SEN net21 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net86 D net25 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX0 net86 c net93 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX5 net94 net93 VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX7 net93 cn net37 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net37 net94 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net94 cn net109 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX19 net53 net118 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net109 c net53 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX21 net118 net109 VDD VNW PHVT11LL_CKT W=0.53u L=40.00n
XX24 SEN SE VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.18u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX23 Q net118 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS SDQV4_12TH40
.SUBCKT SDQV6_12TH40 CK D Q SE SI VDD VSS
XX31 net86 SE net78 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net78 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net82 SEN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX2 net86 D net82 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX3 net86 cn net93 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX4 net94 net93 VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX6 net93 c net102 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net102 net94 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net94 c net109 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX16 net110 net118 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net109 cn net110 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net118 net109 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX25 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX22 Q net118 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX27 net25 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX28 net21 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX29 net86 SEN net21 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net86 D net25 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX0 net86 c net93 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX5 net94 net93 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX7 net93 cn net37 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net37 net94 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net94 cn net109 VNW PHVT11LL_CKT W=0.325u L=40.00n
XX19 net53 net118 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net109 c net53 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX21 net118 net109 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX24 SEN SE VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX23 Q net118 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS SDQV6_12TH40
.SUBCKT SDQV8_12TH40 CK D Q SE SI VDD VSS
XX31 net86 SE net78 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net78 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net82 SEN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX2 net86 D net82 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX3 net86 cn net93 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX4 net94 net93 VSS VPW NHVT11LL_CKT W=0.58u L=40.00n
XX6 net93 c net102 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net102 net94 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net94 c net109 VPW NHVT11LL_CKT W=0.49u L=40.00n
XX16 net110 net118 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net109 cn net110 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net118 net109 VSS VPW NHVT11LL_CKT W=0.66u L=40.00n
XX25 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX22 Q net118 VSS VPW NHVT11LL_CKT W=2.14u L=40.00n
XX27 net25 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX28 net21 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX29 net86 SEN net21 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net86 D net25 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net86 c net93 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX5 net94 net93 VDD VNW PHVT11LL_CKT W=0.49u L=40.00n
XX7 net93 cn net37 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net37 net94 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net94 cn net109 VNW PHVT11LL_CKT W=0.49u L=40.00n
XX19 net53 net118 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net109 c net53 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX21 net118 net109 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX24 SEN SE VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.21u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX23 Q net118 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS SDQV8_12TH40
.SUBCKT SDRNQNV0_12TH40 CK D QN RDN SE SI VDD VSS
XX36 R RDN VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX32 net110 cn net97 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX31 net110 SE net102 VPW NHVT11LL_CKT W=0.14u L=40.00n
XX30 net102 SI VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX0 net106 SEN VSS VPW NHVT11LL_CKT W=0.53u L=40.00n
XX2 net110 D net106 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX25 net122 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX27 net137 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net122 net97 VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX6 net97 c net130 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net130 net122 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net122 c net137 VPW NHVT11LL_CKT W=0.21u L=40.00n
XX16 net138 net140 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net137 cn net138 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net140 net137 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net137 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX35 SEN SE VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX37 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX33 net110 c net97 VNW PHVT11LL_CKT W=0.29u L=40.00n
XX3 net41 SE VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX28 net37 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX29 net110 SEN net37 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net110 D net41 VNW PHVT11LL_CKT W=0.39u L=40.00n
XX26 net69 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX24 net53 R VDD VNW PHVT11LL_CKT W=0.52u L=40.00n
XX5 net122 net97 net53 VNW PHVT11LL_CKT W=0.4u L=40.00n
XX7 net97 cn net57 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net57 net122 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net122 cn net137 VNW PHVT11LL_CKT W=0.24u L=40.00n
XX19 net73 net140 net69 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net137 c net73 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net140 net137 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net137 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=0.18u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.38u L=40.00n
.ENDS SDRNQNV0_12TH40
.SUBCKT SDRNQNV2_12TH40 CK D QN RDN SE SI VDD VSS
XX36 R RDN VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX32 net110 cn net97 VPW NHVT11LL_CKT W=330.00n L=40.00n
XX31 net110 SE net102 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net102 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX0 net106 SEN VSS VPW NHVT11LL_CKT W=0.59u L=40.00n
XX2 net110 D net106 VPW NHVT11LL_CKT W=0.32u L=40.00n
XX25 net122 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX27 net137 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net122 net97 VSS VPW NHVT11LL_CKT W=360.00n L=40.00n
XX6 net97 c net130 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net130 net122 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net122 c net137 VPW NHVT11LL_CKT W=330.00n L=40.00n
XX16 net138 net140 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net137 cn net138 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net140 net137 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net137 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX35 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX37 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX33 net110 c net97 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX3 net41 SE VDD VNW PHVT11LL_CKT W=0.58u L=40.00n
XX28 net37 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX29 net110 SEN net37 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net110 D net41 VNW PHVT11LL_CKT W=0.44u L=40.00n
XX26 net69 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX24 net53 R VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX5 net122 net97 net53 VNW PHVT11LL_CKT W=540.00n L=40.00n
XX7 net97 cn net57 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net57 net122 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net122 cn net137 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX19 net73 net140 net69 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net137 c net73 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net140 net137 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net137 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
.ENDS SDRNQNV2_12TH40
.SUBCKT SDRNQNV4_12TH40 CK D QN RDN SE SI VDD VSS
XX36 R RDN VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX32 net110 cn net97 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX31 net110 SE net102 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net102 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX0 net106 SEN VSS VPW NHVT11LL_CKT W=0.57u L=40.00n
XX2 net110 D net106 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX25 net122 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX27 net137 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net122 net97 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX6 net97 c net130 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net130 net122 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net122 c net137 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX16 net138 net140 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net137 cn net138 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net140 net137 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net137 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX35 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX37 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX33 net110 c net97 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX3 net41 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX28 net37 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX29 net110 SEN net37 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net110 D net41 VNW PHVT11LL_CKT W=0.4u L=40.00n
XX26 net69 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX24 net53 R VDD VNW PHVT11LL_CKT W=0.92u L=40.00n
XX5 net122 net97 net53 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX7 net97 cn net57 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net57 net122 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net122 cn net137 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX19 net73 net140 net69 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net137 c net73 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net140 net137 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net137 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
.ENDS SDRNQNV4_12TH40
.SUBCKT SDRNQNV6_12TH40 CK D QN RDN SE SI VDD VSS
XX36 R RDN VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX32 net110 cn net97 VPW NHVT11LL_CKT W=0.5u L=40.00n
XX31 net110 SE net102 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net102 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX0 net106 SEN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX2 net110 D net106 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX25 net122 R VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX27 net137 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net122 net97 VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX6 net97 c net130 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net130 net122 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net122 c net137 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX16 net138 net140 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net137 cn net138 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net140 net137 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net137 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX35 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX37 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX33 net110 c net97 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX3 net41 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX28 net37 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX29 net110 SEN net37 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net110 D net41 VNW PHVT11LL_CKT W=0.54u L=40.00n
XX26 net69 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX24 net53 R VDD VNW PHVT11LL_CKT W=0.92u L=40.00n
XX5 net122 net97 net53 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX7 net97 cn net57 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net57 net122 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net122 cn net137 VNW PHVT11LL_CKT W=0.52u L=40.00n
XX19 net73 net140 net69 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net137 c net73 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net140 net137 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net137 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
.ENDS SDRNQNV6_12TH40
.SUBCKT SDRNQV0_12TH40 CK D Q RDN SE SI VDD VSS
XX36 R RDN VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX18 net32 net37 VSS VPW NHVT11LL_CKT W=0.185u L=40.00n
XX17 net37 cn net30 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net30 net32 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net46 c net37 VPW NHVT11LL_CKT W=0.21u L=40.00n
XX9 net38 net46 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net77 c net38 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net46 net77 VSS VPW NHVT11LL_CKT W=0.24u L=40.00n
XX27 net37 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net46 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX2 net58 D net62 VPW NHVT11LL_CKT W=0.32u L=40.00n
XX0 net62 SEN VSS VPW NHVT11LL_CKT W=0.42u L=40.00n
XX30 net66 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net58 SE net66 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX32 net58 cn net77 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX35 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 Q net32 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX37 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX21 net32 net37 VDD VNW PHVT11LL_CKT W=0.21u L=40.00n
XX20 net37 c net101 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX19 net101 net32 net105 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX15 net46 cn net37 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX8 net117 net46 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net77 cn net117 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net46 net77 net121 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX24 net121 R VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX26 net105 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX1 net58 D net133 VNW PHVT11LL_CKT W=0.35u L=40.00n
XX29 net58 SEN net137 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX28 net137 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX3 net133 SE VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX33 net58 c net77 VNW PHVT11LL_CKT W=0.25u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.38u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX23 Q net32 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
.ENDS SDRNQV0_12TH40
.SUBCKT SDRNQV2_12TH40 CK D Q RDN SE SI VDD VSS
XX36 R RDN VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX18 net32 net37 VSS VPW NHVT11LL_CKT W=325.00n L=40.00n
XX17 net37 cn net30 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net30 net32 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net46 c net37 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX9 net38 net46 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net77 c net38 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net46 net77 VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX27 net37 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net46 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX2 net58 D net62 VPW NHVT11LL_CKT W=0.35u L=40.00n
XX0 net62 SEN VSS VPW NHVT11LL_CKT W=520.00n L=40.00n
XX30 net66 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net58 SE net66 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX32 net58 cn net77 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX35 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 Q net32 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX37 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX21 net32 net37 VDD VNW PHVT11LL_CKT W=0.355u L=40.00n
XX20 net37 c net101 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX19 net101 net32 net105 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX15 net46 cn net37 VNW PHVT11LL_CKT W=260.00n L=40.00n
XX8 net117 net46 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net77 cn net117 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net46 net77 net121 VNW PHVT11LL_CKT W=460.00n L=40.00n
XX24 net121 R VDD VNW PHVT11LL_CKT W=0.51u L=40.00n
XX26 net105 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX1 net58 D net133 VNW PHVT11LL_CKT W=0.44u L=40.00n
XX29 net58 SEN net137 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX28 net137 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX3 net133 SE VDD VNW PHVT11LL_CKT W=0.58u L=40.00n
XX33 net58 c net77 VNW PHVT11LL_CKT W=0.31u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX23 Q net32 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS SDRNQV2_12TH40
.SUBCKT SDRNQV4_12TH40 CK D Q RDN SE SI VDD VSS
XX36 R RDN VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX18 net32 net37 VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX17 net37 cn net30 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net30 net32 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net46 c net37 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX9 net38 net46 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net77 c net38 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net46 net77 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX27 net37 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net46 R VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX2 net58 D net62 VPW NHVT11LL_CKT W=0.35u L=40.00n
XX0 net62 SEN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX30 net66 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net58 SE net66 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX32 net58 cn net77 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX35 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 Q net32 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX37 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX21 net32 net37 VDD VNW PHVT11LL_CKT W=0.535u L=40.00n
XX20 net37 c net101 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX19 net101 net32 net105 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX15 net46 cn net37 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX8 net117 net46 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net77 cn net117 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net46 net77 net121 VNW PHVT11LL_CKT W=0.425u L=40.00n
XX24 net121 R VDD VNW PHVT11LL_CKT W=0.92u L=40.00n
XX26 net105 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX1 net58 D net133 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX29 net58 SEN net137 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX28 net137 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX3 net133 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX33 net58 c net77 VNW PHVT11LL_CKT W=0.39u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX23 Q net32 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS SDRNQV4_12TH40
.SUBCKT SDRNQV6_12TH40 CK D Q RDN SE SI VDD VSS
XX36 R RDN VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX18 net32 net37 VSS VPW NHVT11LL_CKT W=0.56u L=40.00n
XX17 net37 cn net30 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net30 net32 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net46 c net37 VPW NHVT11LL_CKT W=0.49u L=40.00n
XX9 net38 net46 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net77 c net38 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net46 net77 VSS VPW NHVT11LL_CKT W=0.49u L=40.00n
XX27 net37 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net46 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX2 net58 D net62 VPW NHVT11LL_CKT W=0.34u L=40.00n
XX0 net62 SEN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX30 net66 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net58 SE net66 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX32 net58 cn net77 VPW NHVT11LL_CKT W=0.5u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX35 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 Q net32 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX37 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX21 net32 net37 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX20 net37 c net101 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX19 net101 net32 net105 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX15 net46 cn net37 VNW PHVT11LL_CKT W=0.42u L=40.00n
XX8 net117 net46 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net77 cn net117 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net46 net77 net121 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX24 net121 R VDD VNW PHVT11LL_CKT W=0.92u L=40.00n
XX26 net105 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX1 net58 D net133 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX29 net58 SEN net137 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX28 net137 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX3 net133 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX33 net58 c net77 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX23 Q net32 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS SDRNQV6_12TH40
.SUBCKT SDRNQV8_12TH40 CK D Q RDN SE SI VDD VSS
XX36 R RDN VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX18 net32 net37 VSS VPW NHVT11LL_CKT W=0.72u L=40.00n
XX17 net37 cn net30 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net30 net32 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net46 c net37 VPW NHVT11LL_CKT W=0.49u L=40.00n
XX9 net38 net46 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net77 c net38 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net46 net77 VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX27 net37 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net46 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX2 net58 D net62 VPW NHVT11LL_CKT W=0.37u L=40.00n
XX0 net62 SEN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX30 net66 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net58 SE net66 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX32 net58 cn net77 VPW NHVT11LL_CKT W=0.5u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX35 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 Q net32 VSS VPW NHVT11LL_CKT W=2.14u L=40.00n
XX37 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX21 net32 net37 VDD VNW PHVT11LL_CKT W=0.78u L=40.00n
XX20 net37 c net101 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX19 net101 net32 net105 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX15 net46 cn net37 VNW PHVT11LL_CKT W=0.49u L=40.00n
XX8 net117 net46 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net77 cn net117 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net46 net77 net121 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX24 net121 R VDD VNW PHVT11LL_CKT W=0.92u L=40.00n
XX26 net105 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX1 net58 D net133 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX29 net58 SEN net137 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX28 net137 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX3 net133 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX33 net58 c net77 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.21u L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX23 Q net32 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS SDRNQV8_12TH40
.SUBCKT SDRSNQNV0_12TH40 CK D QN RDN SDN SE SI VDD VSS
XX41 R RDN VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX39 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX1 net102 SE net94 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net94 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 net98 SEN VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX34 net102 D net98 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX32 net106 R VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX31 net153 SDN net106 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 net114 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX27 net130 R net122 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX26 net122 SDN VSS VPW NHVT11LL_CKT W=0.49u L=40.00n
XX3 net102 cn net0140 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX4 net130 net0140 net122 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX6 net0140 c net138 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net138 net130 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX14 net130 c net153 VPW NHVT11LL_CKT W=0.23u L=40.00n
XX16 net154 net156 net114 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net153 cn net154 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX18 net156 net153 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net153 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX42 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX40 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX38 net102 D net13 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX37 net13 SE VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX36 net25 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX35 net102 SEN net25 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX30 net153 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX28 net73 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX25 net49 R VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX24 net130 SDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX0 net102 c net0140 VNW PHVT11LL_CKT W=0.24u L=40.00n
XX5 net130 net0140 net49 VNW PHVT11LL_CKT W=0.365u L=40.00n
XX7 net0140 cn net53 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net53 net130 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.38u L=40.00n
XX15 net130 cn net153 VNW PHVT11LL_CKT W=0.27u L=40.00n
XX19 net77 net156 net73 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net153 c net77 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net156 net153 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net153 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
.ENDS SDRSNQNV0_12TH40
.SUBCKT SDRSNQNV2_12TH40 CK D QN RDN SDN SE SI VDD VSS
XX41 R RDN VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX39 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX1 net102 SE net94 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net94 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 net98 SEN VSS VPW NHVT11LL_CKT W=520.00n L=40.00n
XX34 net102 D net98 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX32 net106 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net153 SDN net106 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 net114 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX27 net130 R net122 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX26 net122 SDN VSS VPW NHVT11LL_CKT W=0.49u L=40.00n
XX3 net102 cn net0140 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX4 net130 net0140 net122 VPW NHVT11LL_CKT W=0.41u L=40.00n
XX6 net0140 c net138 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net138 net130 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX14 net130 c net153 VPW NHVT11LL_CKT W=0.29u L=40.00n
XX16 net154 net156 net114 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net153 cn net154 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX18 net156 net153 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net153 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX42 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX40 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX38 net102 D net13 VNW PHVT11LL_CKT W=0.45u L=40.00n
XX37 net13 SE VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX36 net25 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX35 net102 SEN net25 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX30 net153 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX28 net73 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX25 net49 R VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX24 net130 SDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX0 net102 c net0140 VNW PHVT11LL_CKT W=0.31u L=40.00n
XX5 net130 net0140 net49 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX7 net0140 cn net53 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net53 net130 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX15 net130 cn net153 VNW PHVT11LL_CKT W=0.35u L=40.00n
XX19 net77 net156 net73 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net153 c net77 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net156 net153 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net153 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS SDRSNQNV2_12TH40
.SUBCKT SDRSNQNV4_12TH40 CK D QN RDN SDN SE SI VDD VSS
XX41 R RDN VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX39 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX1 net102 SE net94 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net94 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 net98 SEN VSS VPW NHVT11LL_CKT W=0.58u L=40.00n
XX34 net102 D net98 VPW NHVT11LL_CKT W=0.35u L=40.00n
XX32 net106 R VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX31 net153 SDN net106 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 net114 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX27 net130 R net122 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX26 net122 SDN VSS VPW NHVT11LL_CKT W=0.565u L=40.00n
XX3 net102 cn net0140 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX4 net130 net0140 net122 VPW NHVT11LL_CKT W=0.53u L=40.00n
XX6 net0140 c net138 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net138 net130 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX14 net130 c net153 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX16 net154 net156 net114 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net153 cn net154 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX18 net156 net153 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net153 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX42 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX40 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX38 net102 D net13 VNW PHVT11LL_CKT W=0.6u L=40.00n
XX37 net13 SE VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX36 net25 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX35 net102 SEN net25 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX30 net153 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX28 net73 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX25 net49 R VDD VNW PHVT11LL_CKT W=0.82u L=40.00n
XX24 net130 SDN VDD VNW PHVT11LL_CKT W=0.21u L=40.00n
XX0 net102 c net0140 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX5 net130 net0140 net49 VNW PHVT11LL_CKT W=0.52u L=40.00n
XX7 net0140 cn net53 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net53 net130 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX15 net130 cn net153 VNW PHVT11LL_CKT W=0.41u L=40.00n
XX19 net77 net156 net73 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net153 c net77 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net156 net153 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net153 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS SDRSNQNV4_12TH40
.SUBCKT SDRSNQNV6_12TH40 CK D QN RDN SDN SE SI VDD VSS
XX41 R RDN VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX39 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX1 net102 SE net94 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net94 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 net98 SEN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX34 net102 D net98 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX32 net106 R VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX31 net153 SDN net106 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 net114 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX27 net130 R net122 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX26 net122 SDN VSS VPW NHVT11LL_CKT W=0.48u L=40.00n
XX3 net102 cn net0140 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX4 net130 net0140 net122 VPW NHVT11LL_CKT W=0.5u L=40.00n
XX6 net0140 c net138 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net138 net130 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX14 net130 c net153 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX16 net154 net156 net114 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net153 cn net154 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX18 net156 net153 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net153 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX42 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX40 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX38 net102 D net13 VNW PHVT11LL_CKT W=0.6u L=40.00n
XX37 net13 SE VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX36 net25 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX35 net102 SEN net25 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX30 net153 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX28 net73 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX25 net49 R VDD VNW PHVT11LL_CKT W=0.92u L=40.00n
XX24 net130 SDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX0 net102 c net0140 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX5 net130 net0140 net49 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX7 net0140 cn net53 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net53 net130 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX15 net130 cn net153 VNW PHVT11LL_CKT W=0.53u L=40.00n
XX19 net77 net156 net73 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net153 c net77 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net156 net153 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net153 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS SDRSNQNV6_12TH40
.SUBCKT SDRSNQV0_12TH40 CK D Q RDN SDN SE SI VDD VSS
XX41 R RDN VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX39 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX1 net102 SE net94 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net94 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 net98 SEN VSS VPW NHVT11LL_CKT W=0.6u L=40.00n
XX34 net102 D net98 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX32 net106 R VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX31 net153 SDN net106 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX29 net114 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX27 net130 R net122 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX26 net122 SDN VSS VPW NHVT11LL_CKT W=0.485u L=40.00n
XX3 net102 cn net0139 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX4 net130 net0139 net122 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX6 net0139 c net138 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net138 net130 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX14 net130 c net153 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX16 net154 net156 net114 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net153 cn net154 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX18 net156 net153 VSS VPW NHVT11LL_CKT W=0.175u L=40.00n
XX22 Q net156 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX42 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX40 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX38 net102 D net13 VNW PHVT11LL_CKT W=0.34u L=40.00n
XX37 net13 SE VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX36 net25 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX35 net102 SEN net25 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX30 net153 SDN VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX28 net73 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX25 net49 R VDD VNW PHVT11LL_CKT W=0.525u L=40.00n
XX24 net130 SDN VDD VNW PHVT11LL_CKT W=0.23u L=40.00n
XX0 net102 c net0139 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX5 net130 net0139 net49 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX7 net0139 cn net53 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net53 net130 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.38u L=40.00n
XX15 net130 cn net153 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX19 net77 net156 net73 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net153 c net77 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net156 net153 VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX23 Q net156 VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
.ENDS SDRSNQV0_12TH40
.SUBCKT SDRSNQV2_12TH40 CK D Q RDN SDN SE SI VDD VSS
XX41 R RDN VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX39 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX1 net102 SE net94 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net94 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 net98 SEN VSS VPW NHVT11LL_CKT W=0.6u L=40.00n
XX34 net102 D net98 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX32 net106 R VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX31 net153 SDN net106 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX29 net114 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX27 net130 R net122 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX26 net122 SDN VSS VPW NHVT11LL_CKT W=0.605u L=40.00n
XX3 net102 cn net0139 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX4 net130 net0139 net122 VPW NHVT11LL_CKT W=0.26u L=40.00n
XX6 net0139 c net138 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net138 net130 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=130.00n L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=185.00n L=40.00n
XX14 net130 c net153 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX16 net154 net156 net114 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net153 cn net154 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX18 net156 net153 VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX22 Q net156 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX42 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX40 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX38 net102 D net13 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX37 net13 SE VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX36 net25 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX35 net102 SEN net25 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX30 net153 SDN VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX28 net73 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX25 net49 R VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX24 net130 SDN VDD VNW PHVT11LL_CKT W=0.23u L=40.00n
XX0 net102 c net0139 VNW PHVT11LL_CKT W=260.00n L=40.00n
XX5 net130 net0139 net49 VNW PHVT11LL_CKT W=470.00n L=40.00n
XX7 net0139 cn net53 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net53 net130 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX15 net130 cn net153 VNW PHVT11LL_CKT W=0.32u L=40.00n
XX19 net77 net156 net73 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net153 c net77 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net156 net153 VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX23 Q net156 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS SDRSNQV2_12TH40
.SUBCKT SDRSNQV4_12TH40 CK D Q RDN SDN SE SI VDD VSS
XX41 R RDN VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX39 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX1 net102 SE net94 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net94 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 net98 SEN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX34 net102 D net98 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX32 net106 R VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX31 net153 SDN net106 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX29 net114 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX27 net130 R net122 VPW NHVT11LL_CKT W=0.31u L=40.00n
XX26 net122 SDN VSS VPW NHVT11LL_CKT W=0.605u L=40.00n
XX3 net102 cn net0139 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX4 net130 net0139 net122 VPW NHVT11LL_CKT W=0.31u L=40.00n
XX6 net0139 c net138 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net138 net130 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX14 net130 c net153 VPW NHVT11LL_CKT W=0.31u L=40.00n
XX16 net154 net156 net114 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net153 cn net154 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX18 net156 net153 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX22 Q net156 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX42 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX40 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX38 net102 D net13 VNW PHVT11LL_CKT W=0.53u L=40.00n
XX37 net13 SE VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX36 net25 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX35 net102 SEN net25 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX30 net153 SDN VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX28 net73 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX25 net49 R VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX24 net130 SDN VDD VNW PHVT11LL_CKT W=0.23u L=40.00n
XX0 net102 c net0139 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX5 net130 net0139 net49 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX7 net0139 cn net53 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net53 net130 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.18u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX15 net130 cn net153 VNW PHVT11LL_CKT W=0.37u L=40.00n
XX19 net77 net156 net73 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net153 c net77 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net156 net153 VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX23 Q net156 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS SDRSNQV4_12TH40
.SUBCKT SDRSNQV6_12TH40 CK D Q RDN SDN SE SI VDD VSS
XX41 R RDN VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX39 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX1 net102 SE net94 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net94 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 net98 SEN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX34 net102 D net98 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX32 net106 R VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX31 net153 SDN net106 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX29 net114 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX27 net130 R net122 VPW NHVT11LL_CKT W=0.355u L=40.00n
XX26 net122 SDN VSS VPW NHVT11LL_CKT W=0.605u L=40.00n
XX3 net102 cn net0139 VPW NHVT11LL_CKT W=0.32u L=40.00n
XX4 net130 net0139 net122 VPW NHVT11LL_CKT W=0.355u L=40.00n
XX6 net0139 c net138 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net138 net130 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX14 net130 c net153 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX16 net154 net156 net114 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net153 cn net154 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX18 net156 net153 VSS VPW NHVT11LL_CKT W=0.435u L=40.00n
XX22 Q net156 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX42 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX40 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX38 net102 D net13 VNW PHVT11LL_CKT W=0.6u L=40.00n
XX37 net13 SE VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX36 net25 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX35 net102 SEN net25 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX30 net153 SDN VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX28 net73 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX25 net49 R VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX24 net130 SDN VDD VNW PHVT11LL_CKT W=0.23u L=40.00n
XX0 net102 c net0139 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX5 net130 net0139 net49 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX7 net0139 cn net53 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net53 net130 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX15 net130 cn net153 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX19 net77 net156 net73 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net153 c net77 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net156 net153 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX23 Q net156 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS SDRSNQV6_12TH40
.SUBCKT SDRSNQV8_12TH40 CK D Q RDN SDN SE SI VDD VSS
XX41 R RDN VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX39 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX1 net102 SE net94 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net94 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 net98 SEN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX34 net102 D net98 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX32 net106 R VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX31 net153 SDN net106 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX29 net114 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX27 net130 R net122 VPW NHVT11LL_CKT W=0.355u L=40.00n
XX26 net122 SDN VSS VPW NHVT11LL_CKT W=0.605u L=40.00n
XX3 net102 cn net0139 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX4 net130 net0139 net122 VPW NHVT11LL_CKT W=0.355u L=40.00n
XX6 net0139 c net138 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net138 net130 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX14 net130 c net153 VPW NHVT11LL_CKT W=0.355u L=40.00n
XX16 net154 net156 net114 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net153 cn net154 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX18 net156 net153 VSS VPW NHVT11LL_CKT W=0.64u L=40.00n
XX22 Q net156 VSS VPW NHVT11LL_CKT W=2.14u L=40.00n
XX42 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX40 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX38 net102 D net13 VNW PHVT11LL_CKT W=0.6u L=40.00n
XX37 net13 SE VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX36 net25 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX35 net102 SEN net25 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX30 net153 SDN VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX28 net73 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX25 net49 R VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX24 net130 SDN VDD VNW PHVT11LL_CKT W=0.23u L=40.00n
XX0 net102 c net0139 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX5 net130 net0139 net49 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX7 net0139 cn net53 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net53 net130 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.21u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX15 net130 cn net153 VNW PHVT11LL_CKT W=0.465u L=40.00n
XX19 net77 net156 net73 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net153 c net77 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net156 net153 VDD VNW PHVT11LL_CKT W=0.74u L=40.00n
XX23 Q net156 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS SDRSNQV8_12TH40
.SUBCKT SDSNQNV0_12TH40 CK D QN SDN SE SI VDD VSS
XX4 net94 net0154 net98 VPW NHVT11LL_CKT W=0.31u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX24 net98 SDN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX6 net0154 c net106 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net106 net94 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net94 c net113 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX18 net120 net113 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net113 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX16 net118 net120 net126 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net113 cn net118 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX25 net126 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX35 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net142 SE net134 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net134 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net138 SEN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX3 net142 D net138 VPW NHVT11LL_CKT W=0.31u L=40.00n
XX33 net142 cn net0154 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX5 net94 net0154 VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.38u L=40.00n
XX28 net94 SDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX7 net0154 cn net33 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net33 net94 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net94 cn net113 VNW PHVT11LL_CKT W=0.22u L=40.00n
XX21 net120 net113 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net113 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX29 net113 SDN VDD VNW PHVT11LL_CKT W=0.16u L=40.00n
XX19 net57 net120 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net113 c net57 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX27 net73 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net69 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net142 SEN net69 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX2 net142 D net73 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX32 net142 c net0154 VNW PHVT11LL_CKT W=0.2u L=40.00n
.ENDS SDSNQNV0_12TH40
.SUBCKT SDSNQNV2_12TH40 CK D QN SDN SE SI VDD VSS
XX4 net94 net0154 net98 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=190.00n L=40.00n
XX24 net98 SDN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX6 net0154 c net106 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net106 net94 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net94 c net113 VPW NHVT11LL_CKT W=0.34u L=40.00n
XX18 net120 net113 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net113 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX16 net118 net120 net126 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net113 cn net118 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX25 net126 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX35 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net142 SE net134 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net134 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net138 SEN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX3 net142 D net138 VPW NHVT11LL_CKT W=0.37u L=40.00n
XX33 net142 cn net0154 VPW NHVT11LL_CKT W=330.00n L=40.00n
XX5 net94 net0154 VDD VNW PHVT11LL_CKT W=330.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
XX28 net94 SDN VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX7 net0154 cn net33 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net33 net94 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net94 cn net113 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX21 net120 net113 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net113 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX29 net113 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net57 net120 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net113 c net57 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX27 net73 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net69 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net142 SEN net69 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX2 net142 D net73 VNW PHVT11LL_CKT W=0.44u L=40.00n
XX32 net142 c net0154 VNW PHVT11LL_CKT W=330.00n L=40.00n
.ENDS SDSNQNV2_12TH40
.SUBCKT SDSNQNV4_12TH40 CK D QN SDN SE SI VDD VSS
XX4 net94 net0154 net98 VPW NHVT11LL_CKT W=0.61u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.155u L=40.00n
XX24 net98 SDN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX6 net0154 c net106 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net106 net94 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net94 c net113 VPW NHVT11LL_CKT W=0.39u L=40.00n
XX18 net120 net113 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net113 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX16 net118 net120 net126 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net113 cn net118 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX25 net126 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX35 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net142 SE net134 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net134 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net138 SEN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX3 net142 D net138 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX33 net142 cn net0154 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX5 net94 net0154 VDD VNW PHVT11LL_CKT W=0.38u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX28 net94 SDN VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX7 net0154 cn net33 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net33 net94 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net94 cn net113 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX21 net120 net113 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net113 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX29 net113 SDN VDD VNW PHVT11LL_CKT W=0.16u L=40.00n
XX19 net57 net120 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net113 c net57 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX27 net73 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net69 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net142 SEN net69 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX2 net142 D net73 VNW PHVT11LL_CKT W=0.52u L=40.00n
XX32 net142 c net0154 VNW PHVT11LL_CKT W=0.36u L=40.00n
.ENDS SDSNQNV4_12TH40
.SUBCKT SDSNQNV6_12TH40 CK D QN SDN SE SI VDD VSS
XX4 net94 net0154 net98 VPW NHVT11LL_CKT W=0.61u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX24 net98 SDN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX6 net0154 c net106 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net106 net94 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net94 c net113 VPW NHVT11LL_CKT W=0.49u L=40.00n
XX18 net120 net113 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net113 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX16 net118 net120 net126 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net113 cn net118 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX25 net126 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX35 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net142 SE net134 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net134 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net138 SEN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX3 net142 D net138 VPW NHVT11LL_CKT W=0.42u L=40.00n
XX33 net142 cn net0154 VPW NHVT11LL_CKT W=0.42u L=40.00n
XX5 net94 net0154 VDD VNW PHVT11LL_CKT W=0.51u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.21u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX28 net94 SDN VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX7 net0154 cn net33 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net33 net94 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net94 cn net113 VNW PHVT11LL_CKT W=0.49u L=40.00n
XX21 net120 net113 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net113 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX29 net113 SDN VDD VNW PHVT11LL_CKT W=0.16u L=40.00n
XX19 net57 net120 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net113 c net57 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX27 net73 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net69 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net142 SEN net69 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX2 net142 D net73 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX32 net142 c net0154 VNW PHVT11LL_CKT W=0.5u L=40.00n
.ENDS SDSNQNV6_12TH40
.SUBCKT SDSNQV0_12TH40 CK D Q SDN SE SI VDD VSS
XX33 net10 cn net9 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX31 net10 SE net18 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net18 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net14 SEN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX3 net10 D net14 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX35 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net30 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net53 cn net38 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX16 net38 net40 net30 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX22 Q net40 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX18 net40 net53 VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX14 net74 c net53 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX9 net54 net74 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net9 c net54 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX24 net62 SDN VSS VPW NHVT11LL_CKT W=0.585u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX4 net74 net9 net62 VPW NHVT11LL_CKT W=0.31u L=40.00n
XX27 net85 SE VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX32 net10 c net9 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX0 net89 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net10 SEN net89 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX2 net10 D net85 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX20 net53 c net105 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net105 net40 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX29 net53 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 Q net40 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX21 net40 net53 VDD VNW PHVT11LL_CKT W=0.21u L=40.00n
XX15 net74 cn net53 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX8 net133 net74 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net9 cn net133 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX28 net74 SDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.38u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX5 net74 net9 VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
.ENDS SDSNQV0_12TH40
.SUBCKT SDSNQV2_12TH40 CK D Q SDN SE SI VDD VSS
XX33 net10 cn net9 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX31 net10 SE net18 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net18 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net14 SEN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX3 net10 D net14 VPW NHVT11LL_CKT W=0.29u L=40.00n
XX35 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net30 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net53 cn net38 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX16 net38 net40 net30 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX22 Q net40 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX18 net40 net53 VSS VPW NHVT11LL_CKT W=290.00n L=40.00n
XX14 net74 c net53 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX9 net54 net74 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net9 c net54 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX24 net62 SDN VSS VPW NHVT11LL_CKT W=0.59u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=185.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=130.00n L=40.00n
XX4 net74 net9 net62 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX27 net85 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX32 net10 c net9 VNW PHVT11LL_CKT W=260.00n L=40.00n
XX0 net89 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net10 SEN net89 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX2 net10 D net85 VNW PHVT11LL_CKT W=400.00n L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX20 net53 c net105 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net105 net40 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX29 net53 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 Q net40 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX21 net40 net53 VDD VNW PHVT11LL_CKT W=0.39u L=40.00n
XX15 net74 cn net53 VNW PHVT11LL_CKT W=0.28u L=40.00n
XX8 net133 net74 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net9 cn net133 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX28 net74 SDN VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX5 net74 net9 VDD VNW PHVT11LL_CKT W=0.28u L=40.00n
.ENDS SDSNQV2_12TH40
.SUBCKT SDSNQV4_12TH40 CK D Q SDN SE SI VDD VSS
XX33 net10 cn net9 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX31 net10 SE net18 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net18 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net14 SEN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX3 net10 D net14 VPW NHVT11LL_CKT W=0.32u L=40.00n
XX35 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net30 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net53 cn net38 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX16 net38 net40 net30 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX22 Q net40 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX18 net40 net53 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX14 net74 c net53 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX9 net54 net74 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net9 c net54 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX24 net62 SDN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX4 net74 net9 net62 VPW NHVT11LL_CKT W=0.44u L=40.00n
XX27 net85 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX32 net10 c net9 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX0 net89 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net10 SEN net89 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX2 net10 D net85 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX20 net53 c net105 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net105 net40 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX29 net53 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 Q net40 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX21 net40 net53 VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX15 net74 cn net53 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX8 net133 net74 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net9 cn net133 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX28 net74 SDN VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.18u L=40.00n
XX5 net74 net9 VDD VNW PHVT11LL_CKT W=0.3u L=40.00n
.ENDS SDSNQV4_12TH40
.SUBCKT SDSNQV6_12TH40 CK D Q SDN SE SI VDD VSS
XX33 net10 cn net9 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX31 net10 SE net18 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net18 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net14 SEN VSS VPW NHVT11LL_CKT W=0.6u L=40.00n
XX3 net10 D net14 VPW NHVT11LL_CKT W=0.34u L=40.00n
XX35 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net30 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net53 cn net38 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX16 net38 net40 net30 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX22 Q net40 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX18 net40 net53 VSS VPW NHVT11LL_CKT W=0.44u L=40.00n
XX14 net74 c net53 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX9 net54 net74 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net9 c net54 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX24 net62 SDN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX4 net74 net9 net62 VPW NHVT11LL_CKT W=0.53u L=40.00n
XX27 net85 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX32 net10 c net9 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX0 net89 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net10 SEN net89 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX2 net10 D net85 VNW PHVT11LL_CKT W=0.55u L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX20 net53 c net105 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net105 net40 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX29 net53 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 Q net40 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX21 net40 net53 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX15 net74 cn net53 VNW PHVT11LL_CKT W=0.34u L=40.00n
XX8 net133 net74 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net9 cn net133 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX28 net74 SDN VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX5 net74 net9 VDD VNW PHVT11LL_CKT W=0.37u L=40.00n
.ENDS SDSNQV6_12TH40
.SUBCKT SDSNQV8_12TH40 CK D Q SDN SE SI VDD VSS
XX33 net10 cn net9 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX31 net10 SE net18 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net18 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net14 SEN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX3 net10 D net14 VPW NHVT11LL_CKT W=0.37u L=40.00n
XX35 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net30 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net53 cn net38 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX16 net38 net40 net30 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX22 Q net40 VSS VPW NHVT11LL_CKT W=2.14u L=40.00n
XX18 net40 net53 VSS VPW NHVT11LL_CKT W=0.65u L=40.00n
XX14 net74 c net53 VPW NHVT11LL_CKT W=0.44u L=40.00n
XX9 net54 net74 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net9 c net54 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX24 net62 SDN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX4 net74 net9 net62 VPW NHVT11LL_CKT W=0.61u L=40.00n
XX27 net85 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX32 net10 c net9 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX0 net89 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net10 SEN net89 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX2 net10 D net85 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX20 net53 c net105 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net105 net40 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX29 net53 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 Q net40 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX21 net40 net53 VDD VNW PHVT11LL_CKT W=0.89u L=40.00n
XX15 net74 cn net53 VNW PHVT11LL_CKT W=0.42u L=40.00n
XX8 net133 net74 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net9 cn net133 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX28 net74 SDN VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.21u L=40.00n
XX5 net74 net9 VDD VNW PHVT11LL_CKT W=0.49u L=40.00n
.ENDS SDSNQV8_12TH40
.SUBCKT SDXQNV0_12TH40 CK DA DB QN SA SE SI VDD VSS
XX43 net140 SAN net171 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX6 net103 c net108 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX3 net156 cn net103 VPW NHVT11LL_CKT W=0.29u L=40.00n
XX4 net104 net103 VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX9 net108 net104 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX14 net104 c net123 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX16 net124 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net123 cn net124 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 s net123 VSS VPW NHVT11LL_CKT W=0.17u L=40.00n
XX22 QN s VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX26 net140 DB VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX24 SAN SA VSS VPW NHVT11LL_CKT W=0.255u L=40.00n
XX28 net148 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 net167 SE net148 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX34 net156 net167 VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX32 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX41 net171 SEN net167 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX45 net172 SA net171 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX46 net172 DA VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX0 net156 c net103 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX5 net104 net103 VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX7 net103 cn net19 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net19 net104 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.38u L=40.00n
XX15 net104 cn net123 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX19 net43 s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net123 c net43 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX21 s net123 VDD VNW PHVT11LL_CKT W=0.24u L=40.00n
XX23 QN s VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX44 net140 SA net171 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX25 SAN SA VDD VNW PHVT11LL_CKT W=0.29u L=40.00n
XX27 net140 DB VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX30 net71 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX31 net167 SEN net71 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX33 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX35 net156 net167 VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX42 net171 SE net167 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX47 net172 SAN net171 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX48 net172 DA VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
.ENDS SDXQNV0_12TH40
.SUBCKT SDXQNV2_12TH40 CK DA DB QN SA SE SI VDD VSS
XX43 net140 SAN net171 VPW NHVT11LL_CKT W=150.00n L=40.00n
XX6 net103 c net108 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX3 net156 cn net103 VPW NHVT11LL_CKT W=0.29u L=40.00n
XX4 net104 net103 VSS VPW NHVT11LL_CKT W=355.00n L=40.00n
XX9 net108 net104 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=130.00n L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=185.00n L=40.00n
XX14 net104 c net123 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX16 net124 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net123 cn net124 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 s net123 VSS VPW NHVT11LL_CKT W=0.265u L=40.00n
XX22 QN s VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX26 net140 DB VSS VPW NHVT11LL_CKT W=150.00n L=40.00n
XX24 SAN SA VSS VPW NHVT11LL_CKT W=275.00n L=40.00n
XX28 net148 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 net167 SE net148 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX34 net156 net167 VSS VPW NHVT11LL_CKT W=0.42u L=40.00n
XX32 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX41 net171 SEN net167 VPW NHVT11LL_CKT W=150.00n L=40.00n
XX45 net172 SA net171 VPW NHVT11LL_CKT W=150.00n L=40.00n
XX46 net172 DA VSS VPW NHVT11LL_CKT W=150.00n L=40.00n
XX0 net156 c net103 VNW PHVT11LL_CKT W=260.00n L=40.00n
XX5 net104 net103 VDD VNW PHVT11LL_CKT W=440.00n L=40.00n
XX7 net103 cn net19 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net19 net104 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=130.00n L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX15 net104 cn net123 VNW PHVT11LL_CKT W=260.00n L=40.00n
XX19 net43 s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net123 c net43 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX21 s net123 VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX23 QN s VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX44 net140 SA net171 VNW PHVT11LL_CKT W=260.00n L=40.00n
XX25 SAN SA VDD VNW PHVT11LL_CKT W=315.00n L=40.00n
XX27 net140 DB VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX30 net71 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX31 net167 SEN net71 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX33 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX35 net156 net167 VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
XX42 net171 SE net167 VNW PHVT11LL_CKT W=260.00n L=40.00n
XX47 net172 SAN net171 VNW PHVT11LL_CKT W=260.00n L=40.00n
XX48 net172 DA VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
.ENDS SDXQNV2_12TH40
.SUBCKT SDXQNV4_12TH40 CK DA DB QN SA SE SI VDD VSS
XX43 net140 SAN net171 VPW NHVT11LL_CKT W=0.17u L=40.00n
XX6 net103 c net108 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX3 net156 cn net103 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX4 net104 net103 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX9 net108 net104 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX14 net104 c net123 VPW NHVT11LL_CKT W=0.32u L=40.00n
XX16 net124 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net123 cn net124 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 s net123 VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX22 QN s VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX26 net140 DB VSS VPW NHVT11LL_CKT W=0.17u L=40.00n
XX24 SAN SA VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX28 net148 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 net167 SE net148 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX34 net156 net167 VSS VPW NHVT11LL_CKT W=0.45u L=40.00n
XX32 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX41 net171 SEN net167 VPW NHVT11LL_CKT W=0.17u L=40.00n
XX45 net172 SA net171 VPW NHVT11LL_CKT W=0.17u L=40.00n
XX46 net172 DA VSS VPW NHVT11LL_CKT W=0.17u L=40.00n
XX0 net156 c net103 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX5 net104 net103 VDD VNW PHVT11LL_CKT W=0.52u L=40.00n
XX7 net103 cn net19 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net19 net104 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.18u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX15 net104 cn net123 VNW PHVT11LL_CKT W=0.365u L=40.00n
XX19 net43 s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net123 c net43 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX21 s net123 VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX23 QN s VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX44 net140 SA net171 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX25 SAN SA VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX27 net140 DB VDD VNW PHVT11LL_CKT W=0.55u L=40.00n
XX30 net71 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX31 net167 SEN net71 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX33 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX35 net156 net167 VDD VNW PHVT11LL_CKT W=0.3u L=40.00n
XX42 net171 SE net167 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX47 net172 SAN net171 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX48 net172 DA VDD VNW PHVT11LL_CKT W=0.55u L=40.00n
.ENDS SDXQNV4_12TH40
.SUBCKT SDXQNV6_12TH40 CK DA DB QN SA SE SI VDD VSS
XX43 net140 SAN net171 VPW NHVT11LL_CKT W=0.21u L=40.00n
XX6 net103 c net108 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX3 net156 cn net103 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX4 net104 net103 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX9 net108 net104 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX14 net104 c net123 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX16 net124 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net123 cn net124 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 s net123 VSS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX22 QN s VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX26 net140 DB VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX24 SAN SA VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX28 net148 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 net167 SE net148 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX34 net156 net167 VSS VPW NHVT11LL_CKT W=0.575u L=40.00n
XX32 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX41 net171 SEN net167 VPW NHVT11LL_CKT W=0.21u L=40.00n
XX45 net172 SA net171 VPW NHVT11LL_CKT W=0.21u L=40.00n
XX46 net172 DA VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX0 net156 c net103 VNW PHVT11LL_CKT W=0.33u L=40.00n
XX5 net104 net103 VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX7 net103 cn net19 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net19 net104 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX15 net104 cn net123 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX19 net43 s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net123 c net43 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX21 s net123 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX23 QN s VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX44 net140 SA net171 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX25 SAN SA VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX27 net140 DB VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX30 net71 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX31 net167 SEN net71 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX33 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX35 net156 net167 VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX42 net171 SE net167 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX47 net172 SAN net171 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX48 net172 DA VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
.ENDS SDXQNV6_12TH40
.SUBCKT SDXQV0_12TH40 CK DA DB Q SA SE SI VDD VSS
XX46 net12 DA VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX45 net12 SA net19 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX41 net19 SEN net23 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX32 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX34 net28 net23 VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX29 net23 SE net36 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX28 net36 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX24 SAN SA VSS VPW NHVT11LL_CKT W=0.255u L=40.00n
XX26 net44 DB VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX22 Q net63 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX18 s net63 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net63 cn net56 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net56 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net76 c net63 VPW NHVT11LL_CKT W=0.22u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net72 net76 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net76 net83 VSS VPW NHVT11LL_CKT W=0.34u L=40.00n
XX3 net28 cn net83 VPW NHVT11LL_CKT W=0.29u L=40.00n
XX6 net83 c net72 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX43 net44 SAN net19 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX48 net12 DA VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX47 net12 SAN net19 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX42 net19 SE net23 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX35 net28 net23 VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX33 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX31 net23 SEN net119 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX30 net119 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX27 net44 DB VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX25 SAN SA VDD VNW PHVT11LL_CKT W=0.29u L=40.00n
XX44 net44 SA net19 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX23 Q net63 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX21 s net63 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net63 c net143 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net143 s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net76 cn net63 VNW PHVT11LL_CKT W=0.2u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.38u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net167 net76 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net83 cn net167 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net76 net83 VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX0 net28 c net83 VNW PHVT11LL_CKT W=0.2u L=40.00n
.ENDS SDXQV0_12TH40
.SUBCKT SDXQV2_12TH40 CK DA DB Q SA SE SI VDD VSS
XX46 net12 DA VSS VPW NHVT11LL_CKT W=190.00n L=40.00n
XX45 net12 SA net19 VPW NHVT11LL_CKT W=190.00n L=40.00n
XX41 net19 SEN net23 VPW NHVT11LL_CKT W=190.00n L=40.00n
XX32 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX34 net28 net23 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX29 net23 SE net36 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX28 net36 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX24 SAN SA VSS VPW NHVT11LL_CKT W=300.00n L=40.00n
XX26 net44 DB VSS VPW NHVT11LL_CKT W=190.00n L=40.00n
XX22 Q net63 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX18 s net63 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net63 cn net56 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net56 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net76 c net63 VPW NHVT11LL_CKT W=330.00n L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=190.00n L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net72 net76 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net76 net83 VSS VPW NHVT11LL_CKT W=455.00n L=40.00n
XX3 net28 cn net83 VPW NHVT11LL_CKT W=330.00n L=40.00n
XX6 net83 c net72 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX43 net44 SAN net19 VPW NHVT11LL_CKT W=190.00n L=40.00n
XX48 net12 DA VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX47 net12 SAN net19 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX42 net19 SE net23 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX35 net28 net23 VDD VNW PHVT11LL_CKT W=0.23u L=40.00n
XX33 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX31 net23 SEN net119 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX30 net119 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX27 net44 DB VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX25 SAN SA VDD VNW PHVT11LL_CKT W=340.00n L=40.00n
XX44 net44 SA net19 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX23 Q net63 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX21 s net63 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net63 c net143 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net143 s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net76 cn net63 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net167 net76 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net83 cn net167 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net76 net83 VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX0 net28 c net83 VNW PHVT11LL_CKT W=0.23u L=40.00n
.ENDS SDXQV2_12TH40
.SUBCKT SDXQV4_12TH40 CK DA DB Q SA SE SI VDD VSS
XX46 net12 DA VSS VPW NHVT11LL_CKT W=0.205u L=40.00n
XX45 net12 SA net19 VPW NHVT11LL_CKT W=0.205u L=40.00n
XX41 net19 SEN net23 VPW NHVT11LL_CKT W=0.205u L=40.00n
XX32 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX34 net28 net23 VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX29 net23 SE net36 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX28 net36 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX24 SAN SA VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX26 net44 DB VSS VPW NHVT11LL_CKT W=0.205u L=40.00n
XX22 Q net63 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX18 s net63 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net63 cn net56 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net56 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net76 c net63 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.155u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX9 net72 net76 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net76 net83 VSS VPW NHVT11LL_CKT W=0.46u L=40.00n
XX3 net28 cn net83 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX6 net83 c net72 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX43 net44 SAN net19 VPW NHVT11LL_CKT W=0.205u L=40.00n
XX48 net12 DA VDD VNW PHVT11LL_CKT W=0.55u L=40.00n
XX47 net12 SAN net19 VNW PHVT11LL_CKT W=0.425u L=40.00n
XX42 net19 SE net23 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX35 net28 net23 VDD VNW PHVT11LL_CKT W=0.3u L=40.00n
XX33 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX31 net23 SEN net119 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX30 net119 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX27 net44 DB VDD VNW PHVT11LL_CKT W=0.55u L=40.00n
XX25 SAN SA VDD VNW PHVT11LL_CKT W=0.355u L=40.00n
XX44 net44 SA net19 VNW PHVT11LL_CKT W=0.425u L=40.00n
XX23 Q net63 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX21 s net63 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net63 c net143 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net143 s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net76 cn net63 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX8 net167 net76 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net83 cn net167 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net76 net83 VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX0 net28 c net83 VNW PHVT11LL_CKT W=0.3u L=40.00n
.ENDS SDXQV4_12TH40
.SUBCKT SDXQV6_12TH40 CK DA DB Q SA SE SI VDD VSS
XX46 net12 DA VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX45 net12 SA net19 VPW NHVT11LL_CKT W=0.21u L=40.00n
XX41 net19 SEN net23 VPW NHVT11LL_CKT W=0.21u L=40.00n
XX32 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX34 net28 net23 VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX29 net23 SE net36 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX28 net36 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX24 SAN SA VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX26 net44 DB VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX22 Q net63 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX18 s net63 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net63 cn net56 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net56 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net76 c net63 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX9 net72 net76 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net76 net83 VSS VPW NHVT11LL_CKT W=0.435u L=40.00n
XX3 net28 cn net83 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX6 net83 c net72 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX43 net44 SAN net19 VPW NHVT11LL_CKT W=0.21u L=40.00n
XX48 net12 DA VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX47 net12 SAN net19 VNW PHVT11LL_CKT W=0.44u L=40.00n
XX42 net19 SE net23 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX35 net28 net23 VDD VNW PHVT11LL_CKT W=330.00n L=40.00n
XX33 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX31 net23 SEN net119 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX30 net119 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX27 net44 DB VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX25 SAN SA VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX44 net44 SA net19 VNW PHVT11LL_CKT W=0.44u L=40.00n
XX23 Q net63 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX21 s net63 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net63 c net143 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net143 s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net76 cn net63 VNW PHVT11LL_CKT W=0.44u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.21u L=40.00n
XX8 net167 net76 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net83 cn net167 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net76 net83 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net28 c net83 VNW PHVT11LL_CKT W=330.00n L=40.00n
.ENDS SDXQV6_12TH40
.SUBCKT SDXQV8_12TH40 CK DA DB Q SA SE SI VDD VSS
XX46 net12 DA VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX45 net12 SA net19 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX41 net19 SEN net23 VPW NHVT11LL_CKT W=0.285u L=40.00n
XX32 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX34 net28 net23 VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX29 net23 SE net36 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX28 net36 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX24 SAN SA VSS VPW NHVT11LL_CKT W=0.36u L=40.00n
XX26 net44 DB VSS VPW NHVT11LL_CKT W=0.25u L=40.00n
XX22 Q net63 VSS VPW NHVT11LL_CKT W=2.14u L=40.00n
XX18 s net63 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net63 cn net56 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net56 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net76 c net63 VPW NHVT11LL_CKT W=0.49u L=40.00n
XX12 c cn VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX10 cn CK VSS VPW NHVT11LL_CKT W=0.21u L=40.00n
XX9 net72 net76 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net76 net83 VSS VPW NHVT11LL_CKT W=1u L=40.00n
XX3 net28 cn net83 VPW NHVT11LL_CKT W=0.51u L=40.00n
XX6 net83 c net72 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX43 net44 SAN net19 VPW NHVT11LL_CKT W=0.25u L=40.00n
XX48 net12 DA VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX47 net12 SAN net19 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX42 net19 SE net23 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX35 net28 net23 VDD VNW PHVT11LL_CKT W=0.37u L=40.00n
XX33 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX31 net23 SEN net119 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX30 net119 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX27 net44 DB VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX25 SAN SA VDD VNW PHVT11LL_CKT W=0.415u L=40.00n
XX44 net44 SA net19 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX23 Q net63 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX21 s net63 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net63 c net143 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net143 s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net76 cn net63 VNW PHVT11LL_CKT W=0.49u L=40.00n
XX13 c cn VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX11 cn CK VDD VNW PHVT11LL_CKT W=0.21u L=40.00n
XX8 net167 net76 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net83 cn net167 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net76 net83 VDD VNW PHVT11LL_CKT W=1.21u L=40.00n
XX0 net28 c net83 VNW PHVT11LL_CKT W=0.37u L=40.00n
.ENDS SDXQV8_12TH40
.SUBCKT SEDGRNQNV2_12TH40 CK D E QN RN SE SI VDD VSS
XX10 net227 s net238 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX6 net223 sen VSS VPW NHVT11LL_CKT W=0.52u L=40.00n
XX41 VSS sp net222 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net207 SE net279 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX9 net207 en net227 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX29 VSS m net262 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX28 net262 c pm VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 sen SE VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX35 sp s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX33 m c s VPW NHVT11LL_CKT W=0.33u L=40.00n
XX4 net235 E net238 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX19 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX3 net207 D net235 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX40 net222 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX37 QN s VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX21 net207 cn pm VPW NHVT11LL_CKT W=0.33u L=40.00n
XX23 m pm VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX17 net279 SI VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX13 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX5 net238 RN net223 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX1 net210 en net214 VNW PHVT11LL_CKT W=0.58u L=40.00n
XX2 net207 D net210 VNW PHVT11LL_CKT W=0.58u L=40.00n
XX7 net202 s net214 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX8 net207 E net202 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX0 net214 SE VDD VNW PHVT11LL_CKT W=0.58u L=40.00n
XX11 net207 RN net214 VNW PHVT11LL_CKT W=0.14u L=40.00n
XX14 net186 SI VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net207 sen net186 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net207 c pm VNW PHVT11LL_CKT W=330.00n L=40.00n
XX32 m cn s VNW PHVT11LL_CKT W=0.33u L=40.00n
XX22 m pm VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX34 sp s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX36 QN s VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX12 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX18 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX24 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX30 sen SE VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX26 VDD m net139 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX38 VDD sp net131 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX27 net139 cn pm VNW PHVT11LL_CKT W=120.00n L=40.00n
XX39 net131 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS SEDGRNQNV2_12TH40
.SUBCKT SEDGRNQNV4_12TH40 CK D E QN RN SE SI VDD VSS
XX10 net227 s net238 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX6 net223 sen VSS VPW NHVT11LL_CKT W=0.52u L=40.00n
XX41 VSS sp net222 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net207 SE net279 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX9 net207 en net227 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX29 VSS m net262 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX28 net262 c pm VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 sen SE VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX35 sp s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX33 m c s VPW NHVT11LL_CKT W=0.33u L=40.00n
XX4 net235 E net238 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX19 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX3 net207 D net235 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX40 net222 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX37 QN s VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX21 net207 cn pm VPW NHVT11LL_CKT W=0.33u L=40.00n
XX23 m pm VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX17 net279 SI VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX13 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX5 net238 RN net223 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX1 net210 en net214 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX2 net207 D net210 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX7 net202 s net214 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX8 net207 E net202 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX0 net214 SE VDD VNW PHVT11LL_CKT W=0.585u L=40.00n
XX11 net207 RN net214 VNW PHVT11LL_CKT W=0.14u L=40.00n
XX14 net186 SI VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net207 sen net186 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net207 c pm VNW PHVT11LL_CKT W=330.00n L=40.00n
XX32 m cn s VNW PHVT11LL_CKT W=0.4u L=40.00n
XX22 m pm VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX34 sp s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX36 QN s VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX12 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX18 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX24 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX30 sen SE VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX26 VDD m net139 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX38 VDD sp net131 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX27 net139 cn pm VNW PHVT11LL_CKT W=120.00n L=40.00n
XX39 net131 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS SEDGRNQNV4_12TH40
.SUBCKT SEDGRNQNV6_12TH40 CK D E QN RN SE SI VDD VSS
XX10 net227 s net238 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX6 net223 sen VSS VPW NHVT11LL_CKT W=0.52u L=40.00n
XX41 VSS sp net222 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net207 SE net279 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX9 net207 en net227 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX29 VSS m net262 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX28 net262 c pm VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 sen SE VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX35 sp s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX33 m c s VPW NHVT11LL_CKT W=0.33u L=40.00n
XX4 net235 E net238 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX19 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX3 net207 D net235 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX40 net222 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX37 QN s VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX21 net207 cn pm VPW NHVT11LL_CKT W=0.33u L=40.00n
XX23 m pm VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX17 net279 SI VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX13 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX5 net238 RN net223 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX1 net210 en net214 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX2 net207 D net210 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX7 net202 s net214 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX8 net207 E net202 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX0 net214 SE VDD VNW PHVT11LL_CKT W=0.585u L=40.00n
XX11 net207 RN net214 VNW PHVT11LL_CKT W=0.14u L=40.00n
XX14 net186 SI VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net207 sen net186 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net207 c pm VNW PHVT11LL_CKT W=330.00n L=40.00n
XX32 m cn s VNW PHVT11LL_CKT W=0.48u L=40.00n
XX22 m pm VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX34 sp s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX36 QN s VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX12 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX18 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX24 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX30 sen SE VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX26 VDD m net139 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX38 VDD sp net131 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX27 net139 cn pm VNW PHVT11LL_CKT W=120.00n L=40.00n
XX39 net131 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS SEDGRNQNV6_12TH40
.SUBCKT SEDGRNQV2_12TH40 CK D E Q RN SE SI VDD VSS
XX10 net227 s net238 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX6 net223 sen VSS VPW NHVT11LL_CKT W=0.52u L=40.00n
XX41 VSS sp net222 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net207 SE net279 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX9 net207 en net227 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX29 VSS m net262 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX28 net262 c pm VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 sen SE VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX35 sp s VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX25 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX33 m c s VPW NHVT11LL_CKT W=0.33u L=40.00n
XX4 net235 E net238 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX19 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX3 net207 D net235 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX40 net222 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX37 Q sp VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX21 net207 cn pm VPW NHVT11LL_CKT W=0.33u L=40.00n
XX23 m pm VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX17 net279 SI VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX13 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX5 net238 RN net223 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX1 net210 en net214 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX2 net207 D net210 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX7 net202 s net214 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX8 net207 E net202 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX0 net214 SE VDD VNW PHVT11LL_CKT W=0.585u L=40.00n
XX11 net207 RN net214 VNW PHVT11LL_CKT W=0.14u L=40.00n
XX14 net186 SI VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net207 sen net186 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net207 c pm VNW PHVT11LL_CKT W=330.00n L=40.00n
XX32 m cn s VNW PHVT11LL_CKT W=0.33u L=40.00n
XX22 m pm VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX34 sp s VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX36 Q sp VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX12 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX18 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX24 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX30 sen SE VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX26 VDD m net139 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX38 VDD sp net131 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX27 net139 cn pm VNW PHVT11LL_CKT W=120.00n L=40.00n
XX39 net131 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS SEDGRNQV2_12TH40
.SUBCKT SEDGRNQV4_12TH40 CK D E Q RN SE SI VDD VSS
XX10 net227 s net238 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX6 net223 sen VSS VPW NHVT11LL_CKT W=0.52u L=40.00n
XX41 VSS sp net222 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net207 SE net279 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX9 net207 en net227 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX29 VSS m net262 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX28 net262 c pm VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 sen SE VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX35 sp s VSS VPW NHVT11LL_CKT W=0.36u L=40.00n
XX25 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX33 m c s VPW NHVT11LL_CKT W=0.33u L=40.00n
XX4 net235 E net238 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX19 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX3 net207 D net235 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX40 net222 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX37 Q sp VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX21 net207 cn pm VPW NHVT11LL_CKT W=0.33u L=40.00n
XX23 m pm VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX17 net279 SI VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX13 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX5 net238 RN net223 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX1 net210 en net214 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX2 net207 D net210 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX7 net202 s net214 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX8 net207 E net202 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX0 net214 SE VDD VNW PHVT11LL_CKT W=0.585u L=40.00n
XX11 net207 RN net214 VNW PHVT11LL_CKT W=0.14u L=40.00n
XX14 net186 SI VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net207 sen net186 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net207 c pm VNW PHVT11LL_CKT W=330.00n L=40.00n
XX32 m cn s VNW PHVT11LL_CKT W=0.33u L=40.00n
XX22 m pm VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX34 sp s VDD VNW PHVT11LL_CKT W=0.51u L=40.00n
XX36 Q sp VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX12 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX18 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX24 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX30 sen SE VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX26 VDD m net139 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX38 VDD sp net131 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX27 net139 cn pm VNW PHVT11LL_CKT W=120.00n L=40.00n
XX39 net131 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS SEDGRNQV4_12TH40
.SUBCKT SEDGRNQV6_12TH40 CK D E Q RN SE SI VDD VSS
XX10 net227 s net238 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX6 net223 sen VSS VPW NHVT11LL_CKT W=0.52u L=40.00n
XX41 VSS sp net222 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net207 SE net279 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX9 net207 en net227 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX29 VSS m net262 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX28 net262 c pm VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 sen SE VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX35 sp s VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX25 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX33 m c s VPW NHVT11LL_CKT W=0.33u L=40.00n
XX4 net235 E net238 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX19 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX3 net207 D net235 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX40 net222 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX37 Q sp VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX21 net207 cn pm VPW NHVT11LL_CKT W=0.33u L=40.00n
XX23 m pm VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX17 net279 SI VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX13 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX5 net238 RN net223 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX1 net210 en net214 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX2 net207 D net210 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX7 net202 s net214 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX8 net207 E net202 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX0 net214 SE VDD VNW PHVT11LL_CKT W=0.585u L=40.00n
XX11 net207 RN net214 VNW PHVT11LL_CKT W=0.14u L=40.00n
XX14 net186 SI VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net207 sen net186 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net207 c pm VNW PHVT11LL_CKT W=330.00n L=40.00n
XX32 m cn s VNW PHVT11LL_CKT W=0.33u L=40.00n
XX22 m pm VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX34 sp s VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX36 Q sp VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX12 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX18 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX24 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX30 sen SE VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX26 VDD m net139 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX38 VDD sp net131 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX27 net139 cn pm VNW PHVT11LL_CKT W=120.00n L=40.00n
XX39 net131 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
.ENDS SEDGRNQV6_12TH40
.SUBCKT SEDQNV0_12TH40 CK D E QN SE SI VDD VSS
XX36 VDD ps net188 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX41 net224 c pm VNW PHVT11LL_CKT W=0.33u L=40.00n
XX32 ps s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 net172 cn pm VNW PHVT11LL_CKT W=120.00n L=40.00n
XX22 VDD m net172 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 m pm VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX11 net224 sen net163 VNW PHVT11LL_CKT W=0.12u L=40.00n
XX10 net163 SI VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX6 net224 E net155 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX5 net155 s net143 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX28 m cn s VNW PHVT11LL_CKT W=0.33u L=40.00n
XX37 net188 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
XX3 net224 D net147 VNW PHVT11LL_CKT W=0.59u L=40.00n
XX2 net147 en net143 VNW PHVT11LL_CKT W=0.59u L=40.00n
XX4 net143 SE VDD VNW PHVT11LL_CKT W=0.59u L=40.00n
XX26 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX30 sen SE VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX18 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX16 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX34 QN s VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX29 m c s VPW NHVT11LL_CKT W=0.33u L=40.00n
XX39 VSS ps net271 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX35 QN s VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX38 net271 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 ps s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 VSS m net255 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX24 net255 c pm VPW NHVT11LL_CKT W=120.00n L=40.00n
XX21 m pm VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX9 net231 sen VSS VPW NHVT11LL_CKT W=0.52u L=40.00n
XX40 net224 cn pm VPW NHVT11LL_CKT W=0.33u L=40.00n
XX8 net232 s net231 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX1 net228 E net231 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX0 net224 D net228 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX7 net224 en net232 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX15 net216 SI VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX14 net224 SE net216 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX31 sen SE VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX27 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX19 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX17 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
.ENDS SEDQNV0_12TH40
.SUBCKT SEDQNV2_12TH40 CK D E QN SE SI VDD VSS
XX36 VDD ps net188 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX41 net224 c pm VNW PHVT11LL_CKT W=0.33u L=40.00n
XX32 ps s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 net172 cn pm VNW PHVT11LL_CKT W=120.00n L=40.00n
XX22 VDD m net172 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 m pm VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX11 net224 sen net163 VNW PHVT11LL_CKT W=0.12u L=40.00n
XX10 net163 SI VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX6 net224 E net155 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX5 net155 s net143 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX28 m cn s VNW PHVT11LL_CKT W=0.33u L=40.00n
XX37 net188 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
XX3 net224 D net147 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX2 net147 en net143 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX4 net143 SE VDD VNW PHVT11LL_CKT W=0.585u L=40.00n
XX26 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX30 sen SE VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX18 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX16 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX34 QN s VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX29 m c s VPW NHVT11LL_CKT W=0.33u L=40.00n
XX39 VSS ps net271 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX35 QN s VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX38 net271 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 ps s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 VSS m net255 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX24 net255 c pm VPW NHVT11LL_CKT W=120.00n L=40.00n
XX21 m pm VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX9 net231 sen VSS VPW NHVT11LL_CKT W=0.52u L=40.00n
XX40 net224 cn pm VPW NHVT11LL_CKT W=0.33u L=40.00n
XX8 net232 s net231 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX1 net228 E net231 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX0 net224 D net228 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX7 net224 en net232 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX15 net216 SI VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX14 net224 SE net216 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX31 sen SE VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX27 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX19 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX17 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
.ENDS SEDQNV2_12TH40
.SUBCKT SEDQNV4_12TH40 CK D E QN SE SI VDD VSS
XX36 VDD ps net188 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX41 net224 c pm VNW PHVT11LL_CKT W=0.33u L=40.00n
XX32 ps s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 net172 cn pm VNW PHVT11LL_CKT W=120.00n L=40.00n
XX22 VDD m net172 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 m pm VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX11 net224 sen net163 VNW PHVT11LL_CKT W=0.12u L=40.00n
XX10 net163 SI VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX6 net224 E net155 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX5 net155 s net143 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX28 m cn s VNW PHVT11LL_CKT W=0.42u L=40.00n
XX37 net188 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
XX3 net224 D net147 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX2 net147 en net143 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX4 net143 SE VDD VNW PHVT11LL_CKT W=0.585u L=40.00n
XX26 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX30 sen SE VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX18 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX16 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX34 QN s VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX29 m c s VPW NHVT11LL_CKT W=0.33u L=40.00n
XX39 VSS ps net271 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX35 QN s VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX38 net271 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 ps s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 VSS m net255 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX24 net255 c pm VPW NHVT11LL_CKT W=120.00n L=40.00n
XX21 m pm VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX9 net231 sen VSS VPW NHVT11LL_CKT W=0.52u L=40.00n
XX40 net224 cn pm VPW NHVT11LL_CKT W=0.33u L=40.00n
XX8 net232 s net231 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX1 net228 E net231 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX0 net224 D net228 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX7 net224 en net232 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX15 net216 SI VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX14 net224 SE net216 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX31 sen SE VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX27 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX19 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX17 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
.ENDS SEDQNV4_12TH40
.SUBCKT SEDQNV6_12TH40 CK D E QN SE SI VDD VSS
XX36 VDD ps net188 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX41 net224 c pm VNW PHVT11LL_CKT W=0.33u L=40.00n
XX32 ps s VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 net172 cn pm VNW PHVT11LL_CKT W=120.00n L=40.00n
XX22 VDD m net172 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 m pm VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX11 net224 sen net163 VNW PHVT11LL_CKT W=0.12u L=40.00n
XX10 net163 SI VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX6 net224 E net155 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX5 net155 s net143 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX28 m cn s VNW PHVT11LL_CKT W=0.48u L=40.00n
XX37 net188 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
XX3 net224 D net147 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX2 net147 en net143 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX4 net143 SE VDD VNW PHVT11LL_CKT W=0.585u L=40.00n
XX26 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX30 sen SE VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX18 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX16 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX34 QN s VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX29 m c s VPW NHVT11LL_CKT W=0.33u L=40.00n
XX39 VSS ps net271 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX35 QN s VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX38 net271 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 ps s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 VSS m net255 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX24 net255 c pm VPW NHVT11LL_CKT W=120.00n L=40.00n
XX21 m pm VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX9 net231 sen VSS VPW NHVT11LL_CKT W=0.52u L=40.00n
XX40 net224 cn pm VPW NHVT11LL_CKT W=0.33u L=40.00n
XX8 net232 s net231 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX1 net228 E net231 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX0 net224 D net228 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX7 net224 en net232 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX15 net216 SI VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX14 net224 SE net216 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX31 sen SE VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX27 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX19 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX17 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
.ENDS SEDQNV6_12TH40
.SUBCKT SEDQV0_12TH40 CK D E Q SE SI VDD VSS
XX29 m c s VPW NHVT11LL_CKT W=0.33u L=40.00n
XX39 VSS ps net191 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX35 Q ps VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX38 net191 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 ps s VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX25 VSS m net179 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX24 net179 c pm VPW NHVT11LL_CKT W=120.00n L=40.00n
XX21 m pm VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX9 net155 sen VSS VPW NHVT11LL_CKT W=0.52u L=40.00n
XX40 net148 cn pm VPW NHVT11LL_CKT W=0.33u L=40.00n
XX8 net156 s net155 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX1 net152 E net155 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX0 net148 D net152 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX7 net148 en net156 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX15 net140 SI VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX14 net148 SE net140 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX31 sen SE VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX27 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX19 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX17 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX28 m cn s VNW PHVT11LL_CKT W=0.33u L=40.00n
XX37 net228 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
XX3 net148 D net227 VNW PHVT11LL_CKT W=0.59u L=40.00n
XX2 net227 en net223 VNW PHVT11LL_CKT W=0.59u L=40.00n
XX4 net223 SE VDD VNW PHVT11LL_CKT W=0.59u L=40.00n
XX26 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX30 sen SE VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX18 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX16 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX34 Q ps VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX36 VDD ps net228 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX41 net148 c pm VNW PHVT11LL_CKT W=0.33u L=40.00n
XX32 ps s VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX23 net260 cn pm VNW PHVT11LL_CKT W=120.00n L=40.00n
XX22 VDD m net260 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 m pm VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX11 net148 sen net251 VNW PHVT11LL_CKT W=0.12u L=40.00n
XX10 net251 SI VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX6 net148 E net243 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX5 net243 s net223 VNW PHVT11LL_CKT W=140.00n L=40.00n
.ENDS SEDQV0_12TH40
.SUBCKT SEDQV2_12TH40 CK D E Q SE SI VDD VSS
XX30 sen SE VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX26 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX4 net171 SE VDD VNW PHVT11LL_CKT W=0.585u L=40.00n
XX2 net167 en net171 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX3 net240 D net167 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX37 net160 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
XX28 m cn s VNW PHVT11LL_CKT W=0.33u L=40.00n
XX5 net151 s net171 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX6 net240 E net151 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX10 net143 SI VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX11 net240 sen net143 VNW PHVT11LL_CKT W=0.12u L=40.00n
XX20 m pm VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX22 VDD m net128 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 net128 cn pm VNW PHVT11LL_CKT W=120.00n L=40.00n
XX32 ps s VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX41 net240 c pm VNW PHVT11LL_CKT W=0.33u L=40.00n
XX36 VDD ps net160 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX34 Q ps VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX16 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX18 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX35 Q ps VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX17 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX19 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX27 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX31 sen SE VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX14 net240 SE net248 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX15 net248 SI VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX7 net240 en net232 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX0 net240 D net236 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX1 net236 E net239 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX8 net232 s net239 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX40 net240 cn pm VPW NHVT11LL_CKT W=0.33u L=40.00n
XX9 net239 sen VSS VPW NHVT11LL_CKT W=0.52u L=40.00n
XX21 m pm VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX24 net215 c pm VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 VSS m net215 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 ps s VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX38 net203 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX39 VSS ps net203 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 m c s VPW NHVT11LL_CKT W=0.33u L=40.00n
.ENDS SEDQV2_12TH40
.SUBCKT SEDQV4_12TH40 CK D E Q SE SI VDD VSS
XX30 sen SE VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX26 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX4 net171 SE VDD VNW PHVT11LL_CKT W=0.585u L=40.00n
XX2 net167 en net171 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX3 net240 D net167 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX37 net160 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
XX28 m cn s VNW PHVT11LL_CKT W=0.33u L=40.00n
XX5 net151 s net171 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX6 net240 E net151 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX10 net143 SI VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX11 net240 sen net143 VNW PHVT11LL_CKT W=0.12u L=40.00n
XX20 m pm VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX22 VDD m net128 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 net128 cn pm VNW PHVT11LL_CKT W=120.00n L=40.00n
XX32 ps s VDD VNW PHVT11LL_CKT W=0.51u L=40.00n
XX41 net240 c pm VNW PHVT11LL_CKT W=0.33u L=40.00n
XX36 VDD ps net160 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX34 Q ps VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX16 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX18 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX35 Q ps VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX17 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX19 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX27 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX31 sen SE VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX14 net240 SE net248 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX15 net248 SI VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX7 net240 en net232 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX0 net240 D net236 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX1 net236 E net239 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX8 net232 s net239 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX40 net240 cn pm VPW NHVT11LL_CKT W=0.33u L=40.00n
XX9 net239 sen VSS VPW NHVT11LL_CKT W=0.52u L=40.00n
XX21 m pm VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX24 net215 c pm VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 VSS m net215 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 ps s VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX38 net203 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX39 VSS ps net203 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 m c s VPW NHVT11LL_CKT W=0.33u L=40.00n
.ENDS SEDQV4_12TH40
.SUBCKT SEDQV6_12TH40 CK D E Q SE SI VDD VSS
XX30 sen SE VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX26 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX4 net171 SE VDD VNW PHVT11LL_CKT W=0.585u L=40.00n
XX2 net167 en net171 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX3 net240 D net167 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX37 net160 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
XX28 m cn s VNW PHVT11LL_CKT W=0.33u L=40.00n
XX5 net151 s net171 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX6 net240 E net151 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX10 net143 SI VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX11 net240 sen net143 VNW PHVT11LL_CKT W=0.12u L=40.00n
XX20 m pm VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX22 VDD m net128 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 net128 cn pm VNW PHVT11LL_CKT W=120.00n L=40.00n
XX32 ps s VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX41 net240 c pm VNW PHVT11LL_CKT W=0.33u L=40.00n
XX36 VDD ps net160 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX34 Q ps VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX16 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX18 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX35 Q ps VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX17 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX19 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX27 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX31 sen SE VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX14 net240 SE net248 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX15 net248 SI VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX7 net240 en net232 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX0 net240 D net236 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX1 net236 E net239 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX8 net232 s net239 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX40 net240 cn pm VPW NHVT11LL_CKT W=0.33u L=40.00n
XX9 net239 sen VSS VPW NHVT11LL_CKT W=0.52u L=40.00n
XX21 m pm VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX24 net215 c pm VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 VSS m net215 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 ps s VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX38 net203 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX39 VSS ps net203 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 m c s VPW NHVT11LL_CKT W=0.33u L=40.00n
.ENDS SEDQV6_12TH40
.SUBCKT SEDRNQNV2_12TH40 CK D E QN RDN SE SI VDD VSS
XX46 net176 cn net0485 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX36 ps RDN net104 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX37 net104 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX42 net115 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX43 VSS ps net115 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX32 net124 c s VPW NHVT11LL_CKT W=0.33u L=40.00n
XX39 QN s VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX23 net124 net0485 VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX26 net187 c net0485 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX34 sen SE VSS VPW NHVT11LL_CKT W=0.145u L=40.00n
XX18 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX20 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX16 net148 SI net152 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 net152 RDN VSS VPW NHVT11LL_CKT W=0.52u L=40.00n
XX9 net175 sen net152 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX15 net176 SE net148 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 net176 en net168 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX8 net168 s net175 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX3 net172 E net175 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX2 net176 D net172 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX28 VSS RDN net183 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX27 net183 net124 net187 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX45 net176 c net0485 VNW PHVT11LL_CKT W=0.375u L=40.00n
XX25 net8 cn net0485 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 VDD net124 net8 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX22 net124 net0485 VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX33 sen SE VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX29 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX19 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX17 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX1 net176 D net39 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX0 net39 en net43 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX6 net176 E net47 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX5 net47 s net43 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX21 net0485 RDN VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX12 net176 sen net63 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 net63 SI VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX4 net43 SE VDD VNW PHVT11LL_CKT W=0.585u L=40.00n
XX35 ps s VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX44 ps RDN VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX31 net124 cn s VNW PHVT11LL_CKT W=0.33u L=40.00n
XX40 VDD ps net88 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX41 net88 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
XX38 QN s VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
.ENDS SEDRNQNV2_12TH40
.SUBCKT SEDRNQNV4_12TH40 CK D E QN RDN SE SI VDD VSS
XX46 net176 cn net0485 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX36 ps RDN net104 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX37 net104 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX42 net115 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX43 VSS ps net115 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX32 net124 c s VPW NHVT11LL_CKT W=0.33u L=40.00n
XX39 QN s VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX23 net124 net0485 VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX26 net187 c net0485 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX34 sen SE VSS VPW NHVT11LL_CKT W=0.145u L=40.00n
XX18 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX20 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX16 net148 SI net152 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 net152 RDN VSS VPW NHVT11LL_CKT W=0.52u L=40.00n
XX9 net175 sen net152 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX15 net176 SE net148 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 net176 en net168 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX8 net168 s net175 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX3 net172 E net175 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX2 net176 D net172 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX28 VSS RDN net183 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX27 net183 net124 net187 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX45 net176 c net0485 VNW PHVT11LL_CKT W=0.375u L=40.00n
XX25 net8 cn net0485 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 VDD net124 net8 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX22 net124 net0485 VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX33 sen SE VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX29 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX19 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX17 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX1 net176 D net39 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX0 net39 en net43 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX6 net176 E net47 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX5 net47 s net43 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX21 net0485 RDN VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX12 net176 sen net63 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 net63 SI VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX4 net43 SE VDD VNW PHVT11LL_CKT W=0.585u L=40.00n
XX35 ps s VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX44 ps RDN VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX31 net124 cn s VNW PHVT11LL_CKT W=0.42u L=40.00n
XX40 VDD ps net88 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX41 net88 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
XX38 QN s VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS SEDRNQNV4_12TH40
.SUBCKT SEDRNQNV6_12TH40 CK D E QN RDN SE SI VDD VSS
XX46 net176 cn net0485 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX36 ps RDN net104 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX37 net104 s VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX42 net115 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX43 VSS ps net115 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX32 net124 c s VPW NHVT11LL_CKT W=0.33u L=40.00n
XX39 QN s VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX23 net124 net0485 VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX26 net187 c net0485 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX34 sen SE VSS VPW NHVT11LL_CKT W=0.145u L=40.00n
XX18 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX20 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX16 net148 SI net152 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 net152 RDN VSS VPW NHVT11LL_CKT W=0.52u L=40.00n
XX9 net175 sen net152 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX15 net176 SE net148 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 net176 en net168 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX8 net168 s net175 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX3 net172 E net175 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX2 net176 D net172 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX28 VSS RDN net183 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX27 net183 net124 net187 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX45 net176 c net0485 VNW PHVT11LL_CKT W=0.375u L=40.00n
XX25 net8 cn net0485 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 VDD net124 net8 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX22 net124 net0485 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX33 sen SE VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX29 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX19 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX17 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX1 net176 D net39 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX0 net39 en net43 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX6 net176 E net47 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX5 net47 s net43 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX21 net0485 RDN VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX12 net176 sen net63 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 net63 SI VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX4 net43 SE VDD VNW PHVT11LL_CKT W=0.585u L=40.00n
XX35 ps s VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX44 ps RDN VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX31 net124 cn s VNW PHVT11LL_CKT W=0.48u L=40.00n
XX40 VDD ps net88 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX41 net88 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
XX38 QN s VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS SEDRNQNV6_12TH40
.SUBCKT SEDRNQV2_12TH40 CK D E Q RDN SE SI VDD VSS
XX46 net176 cn net0485 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX36 ps RDN net104 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX37 net104 s VSS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX42 net115 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX43 VSS ps net115 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX32 net124 c s VPW NHVT11LL_CKT W=0.33u L=40.00n
XX39 Q ps VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX23 net124 net0485 VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX26 net187 c net0485 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX34 sen SE VSS VPW NHVT11LL_CKT W=0.145u L=40.00n
XX18 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX20 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX16 net148 SI net152 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 net152 RDN VSS VPW NHVT11LL_CKT W=0.52u L=40.00n
XX9 net175 sen net152 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX15 net176 SE net148 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 net176 en net168 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX8 net168 s net175 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX3 net172 E net175 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX2 net176 D net172 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX28 VSS RDN net183 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX27 net183 net124 net187 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX45 net176 c net0485 VNW PHVT11LL_CKT W=0.375u L=40.00n
XX25 net8 cn net0485 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 VDD net124 net8 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX22 net124 net0485 VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX33 sen SE VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX29 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX19 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX17 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX1 net176 D net39 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX0 net39 en net43 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX6 net176 E net47 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX5 net47 s net43 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX21 net0485 RDN VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX12 net176 sen net63 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 net63 SI VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX4 net43 SE VDD VNW PHVT11LL_CKT W=0.585u L=40.00n
XX35 ps s VDD VNW PHVT11LL_CKT W=0.29u L=40.00n
XX44 ps RDN VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX31 net124 cn s VNW PHVT11LL_CKT W=0.33u L=40.00n
XX40 VDD ps net88 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX41 net88 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
XX38 Q ps VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
.ENDS SEDRNQV2_12TH40
.SUBCKT SEDRNQV4_12TH40 CK D E Q RDN SE SI VDD VSS
XX46 net176 cn net0485 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX36 ps RDN net104 VPW NHVT11LL_CKT W=0.44u L=40.00n
XX37 net104 s VSS VPW NHVT11LL_CKT W=0.44u L=40.00n
XX42 net115 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX43 VSS ps net115 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX32 net124 c s VPW NHVT11LL_CKT W=0.33u L=40.00n
XX39 Q ps VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX23 net124 net0485 VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX26 net187 c net0485 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX34 sen SE VSS VPW NHVT11LL_CKT W=0.145u L=40.00n
XX18 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX20 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX16 net148 SI net152 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 net152 RDN VSS VPW NHVT11LL_CKT W=0.52u L=40.00n
XX9 net175 sen net152 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX15 net176 SE net148 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 net176 en net168 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX8 net168 s net175 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX3 net172 E net175 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX2 net176 D net172 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX28 VSS RDN net183 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX27 net183 net124 net187 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX45 net176 c net0485 VNW PHVT11LL_CKT W=0.375u L=40.00n
XX25 net8 cn net0485 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 VDD net124 net8 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX22 net124 net0485 VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX33 sen SE VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX29 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX19 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX17 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX1 net176 D net39 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX0 net39 en net43 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX6 net176 E net47 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX5 net47 s net43 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX21 net0485 RDN VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX12 net176 sen net63 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 net63 SI VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX4 net43 SE VDD VNW PHVT11LL_CKT W=0.585u L=40.00n
XX35 ps s VDD VNW PHVT11LL_CKT W=0.42u L=40.00n
XX44 ps RDN VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX31 net124 cn s VNW PHVT11LL_CKT W=0.33u L=40.00n
XX40 VDD ps net88 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX41 net88 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
XX38 Q ps VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS SEDRNQV4_12TH40
.SUBCKT SEDRNQV6_12TH40 CK D E Q RDN SE SI VDD VSS
XX46 net176 cn net0485 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX36 ps RDN net104 VPW NHVT11LL_CKT W=0.54u L=40.00n
XX37 net104 s VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX42 net115 cn s VPW NHVT11LL_CKT W=120.00n L=40.00n
XX43 VSS ps net115 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX32 net124 c s VPW NHVT11LL_CKT W=0.33u L=40.00n
XX39 Q ps VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX23 net124 net0485 VSS VPW NHVT11LL_CKT W=0.455u L=40.00n
XX26 net187 c net0485 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 en E VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX34 sen SE VSS VPW NHVT11LL_CKT W=0.145u L=40.00n
XX18 cn CK VSS VPW NHVT11LL_CKT W=0.12u L=40.00n
XX20 c cn VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX16 net148 SI net152 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 net152 RDN VSS VPW NHVT11LL_CKT W=0.52u L=40.00n
XX9 net175 sen net152 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX15 net176 SE net148 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX7 net176 en net168 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX8 net168 s net175 VPW NHVT11LL_CKT W=0.12u L=40.00n
XX3 net172 E net175 VPW NHVT11LL_CKT W=0.52u L=40.00n
XX2 net176 D net172 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX28 VSS RDN net183 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX27 net183 net124 net187 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX45 net176 c net0485 VNW PHVT11LL_CKT W=0.375u L=40.00n
XX25 net8 cn net0485 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX24 VDD net124 net8 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX22 net124 net0485 VDD VNW PHVT11LL_CKT W=0.54u L=40.00n
XX33 sen SE VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX29 en E VDD VNW PHVT11LL_CKT W=0.14u L=40.00n
XX19 c cn VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX17 cn CK VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX1 net176 D net39 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX0 net39 en net43 VNW PHVT11LL_CKT W=0.585u L=40.00n
XX6 net176 E net47 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX5 net47 s net43 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX21 net0485 RDN VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX12 net176 sen net63 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 net63 SI VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX4 net43 SE VDD VNW PHVT11LL_CKT W=0.585u L=40.00n
XX35 ps s VDD VNW PHVT11LL_CKT W=0.49u L=40.00n
XX44 ps RDN VDD VNW PHVT11LL_CKT W=0.12u L=40.00n
XX31 net124 cn s VNW PHVT11LL_CKT W=0.33u L=40.00n
XX40 VDD ps net88 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX41 net88 c s VNW PHVT11LL_CKT W=120.00n L=40.00n
XX38 Q ps VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS SEDRNQV6_12TH40
.SUBCKT SNDQNV2_12TH40 CKN D QN SE SI VDD VSS
XX22 QN net37 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX18 net22 net37 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net37 cn net30 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net30 net22 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net46 c net37 VPW NHVT11LL_CKT W=0.26u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX9 net38 net46 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net53 c net38 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net46 net53 VSS VPW NHVT11LL_CKT W=0.36u L=40.00n
XX3 net54 cn net53 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX2 net54 D net58 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX25 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net58 SEN VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX30 net62 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net54 SE net62 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net37 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX21 net22 net37 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net37 c net93 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net93 net22 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net46 cn net37 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX8 net109 net46 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net53 cn net109 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net46 net53 VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX0 net54 c net53 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX1 net54 D net121 VNW PHVT11LL_CKT W=0.45u L=40.00n
XX29 net54 SEN net125 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX28 net125 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX24 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX27 net121 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
.ENDS SNDQNV2_12TH40
.SUBCKT SNDQNV4_12TH40 CKN D QN SE SI VDD VSS
XX22 QN net37 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX18 net22 net37 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net37 cn net30 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net30 net22 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net46 c net37 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX9 net38 net46 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net53 c net38 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net46 net53 VSS VPW NHVT11LL_CKT W=0.39u L=40.00n
XX3 net54 cn net53 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX2 net54 D net58 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX25 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net58 SEN VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX30 net62 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net54 SE net62 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net37 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX21 net22 net37 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net37 c net93 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net93 net22 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net46 cn net37 VNW PHVT11LL_CKT W=0.415u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX8 net109 net46 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net53 cn net109 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net46 net53 VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX0 net54 c net53 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX1 net54 D net121 VNW PHVT11LL_CKT W=0.52u L=40.00n
XX29 net54 SEN net125 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX28 net125 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX24 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX27 net121 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
.ENDS SNDQNV4_12TH40
.SUBCKT SNDQNV6_12TH40 CKN D QN SE SI VDD VSS
XX22 QN net37 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX18 net22 net37 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net37 cn net30 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net30 net22 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net46 c net37 VPW NHVT11LL_CKT W=330.00n L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX9 net38 net46 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net53 c net38 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net46 net53 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX3 net54 cn net53 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX2 net54 D net58 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX25 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net58 SEN VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX30 net62 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net54 SE net62 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net37 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX21 net22 net37 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net37 c net93 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net93 net22 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net46 cn net37 VNW PHVT11LL_CKT W=0.49u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX8 net109 net46 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net53 cn net109 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net46 net53 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net54 c net53 VNW PHVT11LL_CKT W=0.44u L=40.00n
XX1 net54 D net121 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX29 net54 SEN net125 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX28 net125 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX24 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX27 net121 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
.ENDS SNDQNV6_12TH40
.SUBCKT SNDQV2_12TH40 CKN D Q SE SI VDD VSS
XX31 net94 SE net86 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net86 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net90 SEN VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX25 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net94 D net90 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX3 net94 cn net101 VPW NHVT11LL_CKT W=150.00n L=40.00n
XX4 net102 net101 VSS VPW NHVT11LL_CKT W=360.00n L=40.00n
XX6 net101 c net110 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net110 net102 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX14 net102 c net117 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX16 net118 net126 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net117 cn net118 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net126 net117 VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX22 Q net126 VSS VPW NHVT11LL_CKT W=535.000n L=40.00n
XX27 net33 SE VDD VNW PHVT11LL_CKT W=520.00n L=40.00n
XX24 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX28 net21 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX29 net94 SEN net21 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net94 D net33 VNW PHVT11LL_CKT W=520.00n L=40.00n
XX0 net94 c net101 VNW PHVT11LL_CKT W=260.00n L=40.00n
XX5 net102 net101 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX7 net101 cn net45 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net45 net102 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.4u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX15 net102 cn net117 VNW PHVT11LL_CKT W=260.00n L=40.00n
XX19 net61 net126 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net117 c net61 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX21 net126 net117 VDD VNW PHVT11LL_CKT W=0.29u L=40.00n
XX23 Q net126 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS SNDQV2_12TH40
.SUBCKT SNDQV4_12TH40 CKN D Q SE SI VDD VSS
XX31 net94 SE net86 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net86 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net90 SEN VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX25 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net94 D net90 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX3 net94 cn net101 VPW NHVT11LL_CKT W=0.17u L=40.00n
XX4 net102 net101 VSS VPW NHVT11LL_CKT W=0.39u L=40.00n
XX6 net101 c net110 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net110 net102 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX14 net102 c net117 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX16 net118 net126 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net117 cn net118 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net126 net117 VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX22 Q net126 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX27 net33 SE VDD VNW PHVT11LL_CKT W=0.58u L=40.00n
XX24 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX28 net21 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX29 net94 SEN net21 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net94 D net33 VNW PHVT11LL_CKT W=0.58u L=40.00n
XX0 net94 c net101 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX5 net102 net101 VDD VNW PHVT11LL_CKT W=0.53u L=40.00n
XX7 net101 cn net45 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net45 net102 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.375u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX15 net102 cn net117 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX19 net61 net126 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net117 c net61 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX21 net126 net117 VDD VNW PHVT11LL_CKT W=0.535u L=40.00n
XX23 Q net126 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS SNDQV4_12TH40
.SUBCKT SNDQV6_12TH40 CKN D Q SE SI VDD VSS
XX31 net94 SE net86 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net86 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net90 SEN VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX25 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net94 D net90 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX3 net94 cn net101 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX4 net102 net101 VSS VPW NHVT11LL_CKT W=0.5u L=40.00n
XX6 net101 c net110 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net110 net102 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX14 net102 c net117 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX16 net118 net126 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net117 cn net118 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net126 net117 VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX22 Q net126 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX27 net33 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX24 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX28 net21 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX29 net94 SEN net21 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net94 D net33 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net94 c net101 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX5 net102 net101 VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX7 net101 cn net45 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net45 net102 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX15 net102 cn net117 VNW PHVT11LL_CKT W=0.485u L=40.00n
XX19 net61 net126 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net117 c net61 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX21 net126 net117 VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX23 Q net126 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS SNDQV6_12TH40
.SUBCKT SNDRNQNV2_12TH40 CKN D QN RDN SE SI VDD VSS
XX36 R RDN VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX32 net110 cn net97 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX31 net110 SE net102 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net102 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX0 net106 SEN VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX2 net110 D net106 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX25 net122 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX27 net137 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net122 net97 VSS VPW NHVT11LL_CKT W=360.00n L=40.00n
XX6 net97 c net130 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net130 net122 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net122 c net137 VPW NHVT11LL_CKT W=0.27u L=40.00n
XX16 net138 net140 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net137 cn net138 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net140 net137 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net137 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX35 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX37 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX33 net110 c net97 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX3 net41 SE VDD VNW PHVT11LL_CKT W=0.58u L=40.00n
XX28 net37 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX29 net110 SEN net37 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net110 D net41 VNW PHVT11LL_CKT W=0.44u L=40.00n
XX26 net69 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX24 net53 R VDD VNW PHVT11LL_CKT W=540.00n L=40.00n
XX5 net122 net97 net53 VNW PHVT11LL_CKT W=540.00n L=40.00n
XX7 net97 cn net57 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net57 net122 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net122 cn net137 VNW PHVT11LL_CKT W=330.00n L=40.00n
XX19 net73 net140 net69 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net137 c net73 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net140 net137 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net137 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
.ENDS SNDRNQNV2_12TH40
.SUBCKT SNDRNQNV4_12TH40 CKN D QN RDN SE SI VDD VSS
XX36 R RDN VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX32 net110 cn net97 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX31 net110 SE net102 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net102 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX0 net106 SEN VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX2 net110 D net106 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX25 net122 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX27 net137 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net122 net97 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX6 net97 c net130 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net130 net122 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net122 c net137 VPW NHVT11LL_CKT W=0.28u L=40.00n
XX16 net138 net140 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net137 cn net138 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net140 net137 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net137 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX35 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX37 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX33 net110 c net97 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX3 net41 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX28 net37 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX29 net110 SEN net37 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net110 D net41 VNW PHVT11LL_CKT W=0.49u L=40.00n
XX26 net69 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX24 net53 R VDD VNW PHVT11LL_CKT W=0.92u L=40.00n
XX5 net122 net97 net53 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX7 net97 cn net57 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net57 net122 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net122 cn net137 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX19 net73 net140 net69 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net137 c net73 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net140 net137 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net137 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
.ENDS SNDRNQNV4_12TH40
.SUBCKT SNDRNQNV6_12TH40 CKN D QN RDN SE SI VDD VSS
XX36 R RDN VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX32 net110 cn net97 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX31 net110 SE net102 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net102 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX0 net106 SEN VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX2 net110 D net106 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX25 net122 R VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX27 net137 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net122 net97 VSS VPW NHVT11LL_CKT W=0.42u L=40.00n
XX6 net97 c net130 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net130 net122 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net122 c net137 VPW NHVT11LL_CKT W=330.00n L=40.00n
XX16 net138 net140 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX17 net137 cn net138 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX18 net140 net137 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net137 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX35 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX37 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX33 net110 c net97 VNW PHVT11LL_CKT W=0.44u L=40.00n
XX3 net41 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX28 net37 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX29 net110 SEN net37 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net110 D net41 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX26 net69 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX24 net53 R VDD VNW PHVT11LL_CKT W=0.92u L=40.00n
XX5 net122 net97 net53 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX7 net97 cn net57 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net57 net122 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net122 cn net137 VNW PHVT11LL_CKT W=0.52u L=40.00n
XX19 net73 net140 net69 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net137 c net73 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net140 net137 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net137 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
.ENDS SNDRNQNV6_12TH40
.SUBCKT SNDRNQV2_12TH40 CKN D Q RDN SE SI VDD VSS
XX36 R RDN VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX18 net32 net37 VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX17 net37 cn net30 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net30 net32 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net46 c net37 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX9 net38 net46 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net77 c net38 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net46 net77 VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX27 net37 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net46 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX2 net58 D net62 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX0 net62 SEN VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX30 net66 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net58 SE net66 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX32 net58 cn net77 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=130.00n L=40.00n
XX35 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 Q net32 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX37 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX21 net32 net37 VDD VNW PHVT11LL_CKT W=0.29u L=40.00n
XX20 net37 c net101 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX19 net101 net32 net105 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX15 net46 cn net37 VNW PHVT11LL_CKT W=0.36u L=40.00n
XX8 net117 net46 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net77 cn net117 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net46 net77 net121 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX24 net121 R VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX26 net105 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX1 net58 D net133 VNW PHVT11LL_CKT W=0.44u L=40.00n
XX29 net58 SEN net137 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX28 net137 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX3 net133 SE VDD VNW PHVT11LL_CKT W=0.58u L=40.00n
XX33 net58 c net77 VNW PHVT11LL_CKT W=0.31u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX23 Q net32 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS SNDRNQV2_12TH40
.SUBCKT SNDRNQV4_12TH40 CKN D Q RDN SE SI VDD VSS
XX36 R RDN VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX18 net32 net37 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX17 net37 cn net30 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net30 net32 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net46 c net37 VPW NHVT11LL_CKT W=0.28u L=40.00n
XX9 net38 net46 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net77 c net38 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net46 net77 VSS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX27 net37 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net46 R VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX2 net58 D net62 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX0 net62 SEN VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX30 net66 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net58 SE net66 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX32 net58 cn net77 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX35 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 Q net32 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX37 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX21 net32 net37 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX20 net37 c net101 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX19 net101 net32 net105 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX15 net46 cn net37 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX8 net117 net46 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net77 cn net117 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net46 net77 net121 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX24 net121 R VDD VNW PHVT11LL_CKT W=0.92u L=40.00n
XX26 net105 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX1 net58 D net133 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX29 net58 SEN net137 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX28 net137 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX3 net133 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX33 net58 c net77 VNW PHVT11LL_CKT W=0.37u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX23 Q net32 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS SNDRNQV4_12TH40
.SUBCKT SNDRNQV6_12TH40 CKN D Q RDN SE SI VDD VSS
XX36 R RDN VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX18 net32 net37 VSS VPW NHVT11LL_CKT W=0.56u L=40.00n
XX17 net37 cn net30 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX16 net30 net32 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net46 c net37 VPW NHVT11LL_CKT W=0.32u L=40.00n
XX9 net38 net46 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net77 c net38 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX4 net46 net77 VSS VPW NHVT11LL_CKT W=0.42u L=40.00n
XX27 net37 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net46 R VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX2 net58 D net62 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX0 net62 SEN VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX30 net66 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net58 SE net66 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX32 net58 cn net77 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX35 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 Q net32 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX37 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX21 net32 net37 VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX20 net37 c net101 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX19 net101 net32 net105 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX15 net46 cn net37 VNW PHVT11LL_CKT W=0.42u L=40.00n
XX8 net117 net46 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net77 cn net117 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX5 net46 net77 net121 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX24 net121 R VDD VNW PHVT11LL_CKT W=0.92u L=40.00n
XX26 net105 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX1 net58 D net133 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX29 net58 SEN net137 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX28 net137 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX3 net133 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX33 net58 c net77 VNW PHVT11LL_CKT W=0.43u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX23 Q net32 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS SNDRNQV6_12TH40
.SUBCKT SNDRSNQNV2_12TH40 CKN D QN RDN SDN SE SI VDD VSS
XX41 R RDN VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX39 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX1 net102 SE net94 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net94 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 net98 SEN VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX34 net102 D net98 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX32 net106 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net153 SDN net106 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 net114 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX27 net130 R net122 VPW NHVT11LL_CKT W=0.15u L=40.00n
XX26 net122 SDN VSS VPW NHVT11LL_CKT W=0.49u L=40.00n
XX3 net102 cn net0140 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX4 net130 net0140 net122 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX6 net0140 c net138 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net138 net130 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=130.00n L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX14 net130 c net153 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX16 net154 net156 net114 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net153 cn net154 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX18 net156 net153 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net153 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX42 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX40 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX38 net102 D net13 VNW PHVT11LL_CKT W=0.45u L=40.00n
XX37 net13 SE VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX36 net25 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX35 net102 SEN net25 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX30 net153 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX28 net73 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX25 net49 R VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX24 net130 SDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX0 net102 c net0140 VNW PHVT11LL_CKT W=0.31u L=40.00n
XX5 net130 net0140 net49 VNW PHVT11LL_CKT W=0.49u L=40.00n
XX7 net0140 cn net53 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net53 net130 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX15 net130 cn net153 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX19 net77 net156 net73 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net153 c net77 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net156 net153 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net153 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS SNDRSNQNV2_12TH40
.SUBCKT SNDRSNQNV4_12TH40 CKN D QN RDN SDN SE SI VDD VSS
XX41 R RDN VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX39 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX1 net102 SE net94 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net94 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 net98 SEN VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX34 net102 D net98 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX32 net106 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net153 SDN net106 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 net114 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX27 net130 R net122 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX26 net122 SDN VSS VPW NHVT11LL_CKT W=0.565u L=40.00n
XX3 net102 cn net0140 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX4 net130 net0140 net122 VPW NHVT11LL_CKT W=390.00n L=40.00n
XX6 net0140 c net138 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net138 net130 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX14 net130 c net153 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX16 net154 net156 net114 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net153 cn net154 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX18 net156 net153 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net153 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX42 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX40 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX38 net102 D net13 VNW PHVT11LL_CKT W=0.6u L=40.00n
XX37 net13 SE VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX36 net25 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX35 net102 SEN net25 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX30 net153 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX28 net73 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX25 net49 R VDD VNW PHVT11LL_CKT W=0.82u L=40.00n
XX24 net130 SDN VDD VNW PHVT11LL_CKT W=0.21u L=40.00n
XX0 net102 c net0140 VNW PHVT11LL_CKT W=0.385u L=40.00n
XX5 net130 net0140 net49 VNW PHVT11LL_CKT W=0.57u L=40.00n
XX7 net0140 cn net53 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net53 net130 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX15 net130 cn net153 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX19 net77 net156 net73 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net153 c net77 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net156 net153 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net153 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS SNDRSNQNV4_12TH40
.SUBCKT SNDRSNQNV6_12TH40 CKN D QN RDN SDN SE SI VDD VSS
XX41 R RDN VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX39 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX1 net102 SE net94 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net94 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 net98 SEN VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX34 net102 D net98 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX32 net106 R VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net153 SDN net106 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX29 net114 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX27 net130 R net122 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX26 net122 SDN VSS VPW NHVT11LL_CKT W=0.475u L=40.00n
XX3 net102 cn net0140 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX4 net130 net0140 net122 VPW NHVT11LL_CKT W=0.42u L=40.00n
XX6 net0140 c net138 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net138 net130 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX14 net130 c net153 VPW NHVT11LL_CKT W=0.33u L=40.00n
XX16 net154 net156 net114 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net153 cn net154 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX18 net156 net153 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net153 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX42 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX40 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX38 net102 D net13 VNW PHVT11LL_CKT W=0.6u L=40.00n
XX37 net13 SE VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX36 net25 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX35 net102 SEN net25 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX30 net153 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX28 net73 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX25 net49 R VDD VNW PHVT11LL_CKT W=0.92u L=40.00n
XX24 net130 SDN VDD VNW PHVT11LL_CKT W=0.2u L=40.00n
XX0 net102 c net0140 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX5 net130 net0140 net49 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX7 net0140 cn net53 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net53 net130 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX15 net130 cn net153 VNW PHVT11LL_CKT W=0.53u L=40.00n
XX19 net77 net156 net73 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net153 c net77 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net156 net153 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net153 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS SNDRSNQNV6_12TH40
.SUBCKT SNDRSNQV2_12TH40 CKN D Q RDN SDN SE SI VDD VSS
XX41 R RDN VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX39 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX1 net102 SE net94 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net94 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 net98 SEN VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX34 net102 D net98 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX32 net106 R VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX31 net153 SDN net106 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX29 net114 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX27 net130 R net122 VPW NHVT11LL_CKT W=0.34u L=40.00n
XX26 net122 SDN VSS VPW NHVT11LL_CKT W=0.605u L=40.00n
XX3 net102 cn net0139 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX4 net130 net0139 net122 VPW NHVT11LL_CKT W=0.34u L=40.00n
XX6 net0139 c net138 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net138 net130 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX14 net130 c net153 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX16 net154 net156 net114 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net153 cn net154 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX18 net156 net153 VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX22 Q net156 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX42 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX40 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX38 net102 D net13 VNW PHVT11LL_CKT W=0.44u L=40.00n
XX37 net13 SE VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX36 net25 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX35 net102 SEN net25 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX30 net153 SDN VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX28 net73 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX25 net49 R VDD VNW PHVT11LL_CKT W=0.495u L=40.00n
XX24 net130 SDN VDD VNW PHVT11LL_CKT W=0.245u L=40.00n
XX0 net102 c net0139 VNW PHVT11LL_CKT W=260.00n L=40.00n
XX5 net130 net0139 net49 VNW PHVT11LL_CKT W=0.495u L=40.00n
XX7 net0139 cn net53 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net53 net130 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX15 net130 cn net153 VNW PHVT11LL_CKT W=260.00n L=40.00n
XX19 net77 net156 net73 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net153 c net77 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net156 net153 VDD VNW PHVT11LL_CKT W=0.29u L=40.00n
XX23 Q net156 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS SNDRSNQV2_12TH40
.SUBCKT SNDRSNQV4_12TH40 CKN D Q RDN SDN SE SI VDD VSS
XX41 R RDN VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX39 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX1 net102 SE net94 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net94 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 net98 SEN VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX34 net102 D net98 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX32 net106 R VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX31 net153 SDN net106 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX29 net114 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX27 net130 R net122 VPW NHVT11LL_CKT W=0.385u L=40.00n
XX26 net122 SDN VSS VPW NHVT11LL_CKT W=0.605u L=40.00n
XX3 net102 cn net0139 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX4 net130 net0139 net122 VPW NHVT11LL_CKT W=0.385u L=40.00n
XX6 net0139 c net138 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net138 net130 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.33u L=40.00n
XX14 net130 c net153 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX16 net154 net156 net114 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net153 cn net154 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX18 net156 net153 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX22 Q net156 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX42 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX40 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX38 net102 D net13 VNW PHVT11LL_CKT W=0.53u L=40.00n
XX37 net13 SE VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX36 net25 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX35 net102 SEN net25 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX30 net153 SDN VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX28 net73 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX25 net49 R VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX24 net130 SDN VDD VNW PHVT11LL_CKT W=0.275u L=40.00n
XX0 net102 c net0139 VNW PHVT11LL_CKT W=0.3u L=40.00n
XX5 net130 net0139 net49 VNW PHVT11LL_CKT W=0.56u L=40.00n
XX7 net0139 cn net53 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net53 net130 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX15 net130 cn net153 VNW PHVT11LL_CKT W=0.385u L=40.00n
XX19 net77 net156 net73 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net153 c net77 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net156 net153 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX23 Q net156 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS SNDRSNQV4_12TH40
.SUBCKT SNDRSNQV6_12TH40 CKN D Q RDN SDN SE SI VDD VSS
XX41 R RDN VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX39 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX1 net102 SE net94 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX2 net94 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 net98 SEN VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX34 net102 D net98 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX32 net106 R VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX31 net153 SDN net106 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX29 net114 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX27 net130 R net122 VPW NHVT11LL_CKT W=0.42u L=40.00n
XX26 net122 SDN VSS VPW NHVT11LL_CKT W=0.605u L=40.00n
XX3 net102 cn net0139 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX4 net130 net0139 net122 VPW NHVT11LL_CKT W=0.42u L=40.00n
XX6 net0139 c net138 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net138 net130 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX14 net130 c net153 VPW NHVT11LL_CKT W=0.32u L=40.00n
XX16 net154 net156 net114 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net153 cn net154 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX18 net156 net153 VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX22 Q net156 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX42 R RDN VDD VNW PHVT11LL_CKT W=250.00n L=40.00n
XX40 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX38 net102 D net13 VNW PHVT11LL_CKT W=0.6u L=40.00n
XX37 net13 SE VDD VNW PHVT11LL_CKT W=0.6u L=40.00n
XX36 net25 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX35 net102 SEN net25 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX30 net153 SDN VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX28 net73 R VDD VNW PHVT11LL_CKT W=160.00n L=40.00n
XX25 net49 R VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX24 net130 SDN VDD VNW PHVT11LL_CKT W=0.25u L=40.00n
XX0 net102 c net0139 VNW PHVT11LL_CKT W=0.38u L=40.00n
XX5 net130 net0139 net49 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX7 net0139 cn net53 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net53 net130 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX15 net130 cn net153 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX19 net77 net156 net73 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX20 net153 c net77 VNW PHVT11LL_CKT W=160.00n L=40.00n
XX21 net156 net153 VDD VNW PHVT11LL_CKT W=0.545u L=40.00n
XX23 Q net156 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS SNDRSNQV6_12TH40
.SUBCKT SNDSNQNV2_12TH40 CKN D QN SDN SE SI VDD VSS
XX4 net94 net0154 net98 VPW NHVT11LL_CKT W=0.36u L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX24 net98 SDN VSS VPW NHVT11LL_CKT W=510.00n L=40.00n
XX6 net0154 c net106 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net106 net94 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net94 c net113 VPW NHVT11LL_CKT W=0.26u L=40.00n
XX18 net120 net113 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net113 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX16 net118 net120 net126 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net113 cn net118 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX25 net126 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX35 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net142 SE net134 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net134 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net138 SEN VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX3 net142 D net138 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX33 net142 cn net0154 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX5 net94 net0154 VDD VNW PHVT11LL_CKT W=0.455u L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX28 net94 SDN VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX7 net0154 cn net33 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net33 net94 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net94 cn net113 VNW PHVT11LL_CKT W=0.375u L=40.00n
XX21 net120 net113 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net113 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX29 net113 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net57 net120 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net113 c net57 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX27 net73 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net69 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net142 SEN net69 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX2 net142 D net73 VNW PHVT11LL_CKT W=360.00n L=40.00n
XX32 net142 c net0154 VNW PHVT11LL_CKT W=330.00n L=40.00n
.ENDS SNDSNQNV2_12TH40
.SUBCKT SNDSNQNV4_12TH40 CKN D QN SDN SE SI VDD VSS
XX4 net94 net0154 net98 VPW NHVT11LL_CKT W=0.39u L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX24 net98 SDN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX6 net0154 c net106 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net106 net94 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net94 c net113 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX18 net120 net113 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net113 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX16 net118 net120 net126 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net113 cn net118 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX25 net126 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX35 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net142 SE net134 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net134 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net138 SEN VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX3 net142 D net138 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX33 net142 cn net0154 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX5 net94 net0154 VDD VNW PHVT11LL_CKT W=0.51u L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX28 net94 SDN VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX7 net0154 cn net33 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net33 net94 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net94 cn net113 VNW PHVT11LL_CKT W=0.415u L=40.00n
XX21 net120 net113 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net113 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX29 net113 SDN VDD VNW PHVT11LL_CKT W=0.16u L=40.00n
XX19 net57 net120 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net113 c net57 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX27 net73 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net69 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net142 SEN net69 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX2 net142 D net73 VNW PHVT11LL_CKT W=0.48u L=40.00n
XX32 net142 c net0154 VNW PHVT11LL_CKT W=0.36u L=40.00n
.ENDS SNDSNQNV4_12TH40
.SUBCKT SNDSNQNV6_12TH40 CKN D QN SDN SE SI VDD VSS
XX4 net94 net0154 net98 VPW NHVT11LL_CKT W=0.43u L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.35u L=40.00n
XX24 net98 SDN VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX6 net0154 c net106 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 net106 net94 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX14 net94 c net113 VPW NHVT11LL_CKT W=330.00n L=40.00n
XX18 net120 net113 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX22 QN net113 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX16 net118 net120 net126 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net113 cn net118 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX25 net126 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX35 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net142 SE net134 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX30 net134 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX26 net138 SEN VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX3 net142 D net138 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX33 net142 cn net0154 VPW NHVT11LL_CKT W=0.18u L=40.00n
XX5 net94 net0154 VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX28 net94 SDN VDD VNW PHVT11LL_CKT W=0.22u L=40.00n
XX7 net0154 cn net33 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX8 net33 net94 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX15 net94 cn net113 VNW PHVT11LL_CKT W=0.49u L=40.00n
XX21 net120 net113 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 QN net113 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX29 net113 SDN VDD VNW PHVT11LL_CKT W=0.16u L=40.00n
XX19 net57 net120 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX20 net113 c net57 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX27 net73 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX0 net69 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX1 net142 SEN net69 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX2 net142 D net73 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX32 net142 c net0154 VNW PHVT11LL_CKT W=0.5u L=40.00n
.ENDS SNDSNQNV6_12TH40
.SUBCKT SNDSNQV2_12TH40 CKN D Q SDN SE SI VDD VSS
XX35 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 net22 D net18 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX32 net18 SEN VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX30 net14 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net22 SE net14 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net34 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net57 cn net42 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX16 net42 net44 net34 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX22 Q net44 VSS VPW NHVT11LL_CKT W=535.00n L=40.00n
XX18 net44 net57 VSS VPW NHVT11LL_CKT W=325.00n L=40.00n
XX14 net70 c net57 VPW NHVT11LL_CKT W=260.00n L=40.00n
XX9 net58 net70 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net77 c net58 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX24 net66 net77 VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.3u L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX4 net70 SDN net66 VPW NHVT11LL_CKT W=400.00n L=40.00n
XX3 net22 cn net77 VPW NHVT11LL_CKT W=150.00n L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX26 net85 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX2 net22 D net97 VNW PHVT11LL_CKT W=0.53u L=40.00n
XX1 net97 SE VDD VNW PHVT11LL_CKT W=0.53u L=40.00n
XX27 net22 SEN net85 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX20 net57 c net109 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net109 net44 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX29 net57 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 Q net44 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX21 net44 net57 VDD VNW PHVT11LL_CKT W=325.00n L=40.00n
XX15 net70 cn net57 VNW PHVT11LL_CKT W=260.00n L=40.00n
XX8 net137 net70 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net77 cn net137 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX28 net70 SDN VDD VNW PHVT11LL_CKT W=260.00n L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=350.00n L=40.00n
XX5 net70 net77 VDD VNW PHVT11LL_CKT W=0.36u L=40.00n
XX0 net22 c net77 VNW PHVT11LL_CKT W=260.00n L=40.00n
.ENDS SNDSNQV2_12TH40
.SUBCKT SNDSNQV4_12TH40 CKN D Q SDN SE SI VDD VSS
XX35 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 net22 D net18 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX32 net18 SEN VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX30 net14 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net22 SE net14 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net34 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net57 cn net42 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX16 net42 net44 net34 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX22 Q net44 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX18 net44 net57 VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX14 net70 c net57 VPW NHVT11LL_CKT W=0.3u L=40.00n
XX9 net58 net70 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net77 c net58 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX24 net66 net77 VSS VPW NHVT11LL_CKT W=0.46u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.14u L=40.00n
XX4 net70 SDN net66 VPW NHVT11LL_CKT W=0.46u L=40.00n
XX3 net22 cn net77 VPW NHVT11LL_CKT W=0.17u L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX26 net85 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX2 net22 D net97 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX1 net97 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX27 net22 SEN net85 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX20 net57 c net109 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net109 net44 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX29 net57 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 Q net44 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX21 net44 net57 VDD VNW PHVT11LL_CKT W=0.535u L=40.00n
XX15 net70 cn net57 VNW PHVT11LL_CKT W=0.35u L=40.00n
XX8 net137 net70 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net77 cn net137 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX28 net70 SDN VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.375u L=40.00n
XX5 net70 net77 VDD VNW PHVT11LL_CKT W=0.48u L=40.00n
XX0 net22 c net77 VNW PHVT11LL_CKT W=0.3u L=40.00n
.ENDS SNDSNQV4_12TH40
.SUBCKT SNDSNQV6_12TH40 CKN D Q SDN SE SI VDD VSS
XX35 SEN SE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX33 net22 D net18 VPW NHVT11LL_CKT W=0.2u L=40.00n
XX32 net18 SEN VSS VPW NHVT11LL_CKT W=0.2u L=40.00n
XX30 net14 SI VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX31 net22 SE net14 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX25 net34 SDN VSS VPW NHVT11LL_CKT W=160.00n L=40.00n
XX17 net57 cn net42 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX16 net42 net44 net34 VPW NHVT11LL_CKT W=160.00n L=40.00n
XX22 Q net44 VSS VPW NHVT11LL_CKT W=1.605u L=40.00n
XX18 net44 net57 VSS VPW NHVT11LL_CKT W=0.56u L=40.00n
XX14 net70 c net57 VPW NHVT11LL_CKT W=0.38u L=40.00n
XX9 net58 net70 VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX6 net77 c net58 VPW NHVT11LL_CKT W=120.00n L=40.00n
XX24 net66 net77 VSS VPW NHVT11LL_CKT W=0.57u L=40.00n
XX12 cn c VSS VPW NHVT11LL_CKT W=0.32u L=40.00n
XX10 c CKN VSS VPW NHVT11LL_CKT W=0.15u L=40.00n
XX4 net70 SDN net66 VPW NHVT11LL_CKT W=0.57u L=40.00n
XX3 net22 cn net77 VPW NHVT11LL_CKT W=0.21u L=40.00n
XX34 SEN SE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX26 net85 SI VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
XX2 net22 D net97 VNW PHVT11LL_CKT W=0.61u L=40.00n
XX1 net97 SE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX27 net22 SEN net85 VNW PHVT11LL_CKT W=140.00n L=40.00n
XX20 net57 c net109 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX19 net109 net44 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX29 net57 SDN VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX23 Q net44 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX21 net44 net57 VDD VNW PHVT11LL_CKT W=0.56u L=40.00n
XX15 net70 cn net57 VNW PHVT11LL_CKT W=0.445u L=40.00n
XX8 net137 net70 VDD VNW PHVT11LL_CKT W=120.00n L=40.00n
XX7 net77 cn net137 VNW PHVT11LL_CKT W=120.00n L=40.00n
XX28 net70 SDN VDD VNW PHVT11LL_CKT W=0.445u L=40.00n
XX13 cn c VDD VNW PHVT11LL_CKT W=0.15u L=40.00n
XX11 c CKN VDD VNW PHVT11LL_CKT W=0.425u L=40.00n
XX5 net70 net77 VDD VNW PHVT11LL_CKT W=0.545u L=40.00n
XX0 net22 c net77 VNW PHVT11LL_CKT W=0.38u L=40.00n
.ENDS SNDSNQV6_12TH40
.SUBCKT TBUFV12_12TH40 I OE Z VDD VSS
XX8 Z net034 VSS VPW NHVT11LL_CKT W=3.21u L=40.00n
XX7 net034 OEN VSS VPW NHVT11LL_CKT W=0.8u L=40.00n
XX5 net034 I VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX2 net061 OE net034 VPW NHVT11LL_CKT W=0.8u L=40.00n
XX1 OEN OE VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX9 Z net061 VDD VNW PHVT11LL_CKT W=3.03u L=40.00n
XX6 net061 OE VDD VNW PHVT11LL_CKT W=0.92u L=40.00n
XX4 net061 I VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX3 net034 OEN net061 VNW PHVT11LL_CKT W=0.92u L=40.00n
XX0 OEN OE VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
.ENDS TBUFV12_12TH40
.SUBCKT TBUFV16_12TH40 I OE Z VDD VSS
XX8 Z net034 VSS VPW NHVT11LL_CKT W=3.76u L=40.00n
XX7 net034 OEN VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX5 net034 I VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX2 net061 OE net034 VPW NHVT11LL_CKT W=1.07u L=40.00n
XX1 OEN OE VSS VPW NHVT11LL_CKT W=0.72u L=40.00n
XX9 Z net061 VDD VNW PHVT11LL_CKT W=4.04u L=40.00n
XX6 net061 OE VDD VNW PHVT11LL_CKT W=1.01u L=40.00n
XX4 net061 I VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX3 net034 OEN net061 VNW PHVT11LL_CKT W=1.01u L=40.00n
XX0 OEN OE VDD VNW PHVT11LL_CKT W=0.81u L=40.00n
.ENDS TBUFV16_12TH40
.SUBCKT TBUFV20_12TH40 I OE Z VDD VSS
XX8 Z net034 VSS VPW NHVT11LL_CKT W=4.5u L=40.00n
XX7 net034 OEN VSS VPW NHVT11LL_CKT W=1.47u L=40.00n
XX5 net034 I VSS VPW NHVT11LL_CKT W=2.7u L=40.00n
XX2 net061 OE net034 VPW NHVT11LL_CKT W=1.47u L=40.00n
XX1 OEN OE VSS VPW NHVT11LL_CKT W=0.96u L=40.00n
XX9 Z net061 VDD VNW PHVT11LL_CKT W=5.05u L=40.00n
XX6 net061 OE VDD VNW PHVT11LL_CKT W=1.515u L=40.00n
XX4 net061 I VDD VNW PHVT11LL_CKT W=3.36u L=40.00n
XX3 net034 OEN net061 VNW PHVT11LL_CKT W=1.59u L=40.00n
XX0 OEN OE VDD VNW PHVT11LL_CKT W=1.12u L=40.00n
.ENDS TBUFV20_12TH40
.SUBCKT TBUFV24_12TH40 I OE Z VDD VSS
XX8 Z net034 VSS VPW NHVT11LL_CKT W=5.4u L=40.00n
XX7 net034 OEN VSS VPW NHVT11LL_CKT W=1.47u L=40.00n
XX5 net034 I VSS VPW NHVT11LL_CKT W=2.7u L=40.00n
XX2 net061 OE net034 VPW NHVT11LL_CKT W=1.47u L=40.00n
XX1 OEN OE VSS VPW NHVT11LL_CKT W=0.96u L=40.00n
XX9 Z net061 VDD VNW PHVT11LL_CKT W=6.06u L=40.00n
XX6 net061 OE VDD VNW PHVT11LL_CKT W=1.515u L=40.00n
XX4 net061 I VDD VNW PHVT11LL_CKT W=3.36u L=40.00n
XX3 net034 OEN net061 VNW PHVT11LL_CKT W=1.59u L=40.00n
XX0 OEN OE VDD VNW PHVT11LL_CKT W=1.12u L=40.00n
.ENDS TBUFV24_12TH40
.SUBCKT TBUFV2_12TH40 I OE Z VDD VSS
XX8 Z net034 VSS VPW NHVT11LL_CKT W=530.00n L=40.00n
XX7 net034 OEN VSS VPW NHVT11LL_CKT W=135.00n L=40.00n
XX5 net034 I VSS VPW NHVT11LL_CKT W=270.00n L=40.00n
XX2 net061 OE net034 VPW NHVT11LL_CKT W=135.00n L=40.00n
XX1 OEN OE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 Z net061 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX6 net061 OE VDD VNW PHVT11LL_CKT W=155.00n L=40.00n
XX4 net061 I VDD VNW PHVT11LL_CKT W=305.00n L=40.00n
XX3 net034 OEN net061 VNW PHVT11LL_CKT W=155.00n L=40.00n
XX0 OEN OE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
.ENDS TBUFV2_12TH40
.SUBCKT TBUFV32_12TH40 I OE Z VDD VSS
XX8 Z net034 VSS VPW NHVT11LL_CKT W=7.52u L=40.00n
XX7 net034 OEN VSS VPW NHVT11LL_CKT W=2.14u L=40.00n
XX5 net034 I VSS VPW NHVT11LL_CKT W=4.32u L=40.00n
XX2 net061 OE net034 VPW NHVT11LL_CKT W=2.14u L=40.00n
XX1 OEN OE VSS VPW NHVT11LL_CKT W=1.41u L=40.00n
XX9 Z net061 VDD VNW PHVT11LL_CKT W=8.08u L=40.00n
XX6 net061 OE VDD VNW PHVT11LL_CKT W=2.02u L=40.00n
XX4 net061 I VDD VNW PHVT11LL_CKT W=4.88u L=40.00n
XX3 net034 OEN net061 VNW PHVT11LL_CKT W=2.02u L=40.00n
XX0 OEN OE VDD VNW PHVT11LL_CKT W=1.62u L=40.00n
.ENDS TBUFV32_12TH40
.SUBCKT TBUFV3_12TH40 I OE Z VDD VSS
XX8 Z net034 VSS VPW NHVT11LL_CKT W=0.75u L=40.00n
XX7 net034 OEN VSS VPW NHVT11LL_CKT W=0.19u L=40.00n
XX5 net034 I VSS VPW NHVT11LL_CKT W=0.375u L=40.00n
XX2 net061 OE net034 VPW NHVT11LL_CKT W=0.19u L=40.00n
XX1 OEN OE VSS VPW NHVT11LL_CKT W=120.00n L=40.00n
XX9 Z net061 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX6 net061 OE VDD VNW PHVT11LL_CKT W=0.215u L=40.00n
XX4 net061 I VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX3 net034 OEN net061 VNW PHVT11LL_CKT W=0.215u L=40.00n
XX0 OEN OE VDD VNW PHVT11LL_CKT W=140.00n L=40.00n
.ENDS TBUFV3_12TH40
.SUBCKT TBUFV4_12TH40 I OE Z VDD VSS
XX8 Z net034 VSS VPW NHVT11LL_CKT W=0.94u L=40.00n
XX7 net034 OEN VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX5 net034 I VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX2 net061 OE net034 VPW NHVT11LL_CKT W=0.27u L=40.00n
XX1 OEN OE VSS VPW NHVT11LL_CKT W=0.18u L=40.00n
XX9 Z net061 VDD VNW PHVT11LL_CKT W=1.14u L=40.00n
XX6 net061 OE VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX4 net061 I VDD VNW PHVT11LL_CKT W=0.61u L=40.00n
XX3 net034 OEN net061 VNW PHVT11LL_CKT W=0.305u L=40.00n
XX0 OEN OE VDD VNW PHVT11LL_CKT W=0.205u L=40.00n
.ENDS TBUFV4_12TH40
.SUBCKT TBUFV6_12TH40 I OE Z VDD VSS
XX8 Z net034 VSS VPW NHVT11LL_CKT W=1.41u L=40.00n
XX7 net034 OEN VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX5 net034 I VSS VPW NHVT11LL_CKT W=0.8u L=40.00n
XX2 net061 OE net034 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX1 OEN OE VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX9 Z net061 VDD VNW PHVT11LL_CKT W=1.71u L=40.00n
XX6 net061 OE VDD VNW PHVT11LL_CKT W=0.46u L=40.00n
XX4 net061 I VDD VNW PHVT11LL_CKT W=0.92u L=40.00n
XX3 net034 OEN net061 VNW PHVT11LL_CKT W=0.46u L=40.00n
XX0 OEN OE VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
.ENDS TBUFV6_12TH40
.SUBCKT TBUFV8_12TH40 I OE Z VDD VSS
XX8 Z net034 VSS VPW NHVT11LL_CKT W=1.88u L=40.00n
XX7 net034 OEN VSS VPW NHVT11LL_CKT W=0.535u L=40.00n
XX5 net034 I VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX2 net061 OE net034 VPW NHVT11LL_CKT W=0.535u L=40.00n
XX1 OEN OE VSS VPW NHVT11LL_CKT W=0.355u L=40.00n
XX9 Z net061 VDD VNW PHVT11LL_CKT W=2.28u L=40.00n
XX6 net061 OE VDD VNW PHVT11LL_CKT W=0.505u L=40.00n
XX4 net061 I VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX3 net034 OEN net061 VNW PHVT11LL_CKT W=0.505u L=40.00n
XX0 OEN OE VDD VNW PHVT11LL_CKT W=0.41u L=40.00n
.ENDS TBUFV8_12TH40
.SUBCKT XNOR2V0_12TH40 A1 A2 ZN VDD VSS
XX7 net36 A1N ZN VPW NHVT11LL_CKT W=0.25u L=40.00n
XX6 net24 A1 ZN VPW NHVT11LL_CKT W=0.25u L=40.00n
XX2 net36 A2 VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX0 A1N A1 VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX5 net24 net36 VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX8 net24 A1N ZN VNW PHVT11LL_CKT W=0.25u L=40.00n
XX9 net36 A1 ZN VNW PHVT11LL_CKT W=0.25u L=40.00n
XX3 A1N A1 VDD VNW PHVT11LL_CKT W=0.26u L=40.00n
XX1 net36 A2 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX4 net24 net36 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
.ENDS XNOR2V0_12TH40
.SUBCKT XNOR2V1_12TH40 A1 A2 ZN VDD VSS
XX7 net36 A1N ZN VPW NHVT11LL_CKT W=0.35u L=40.00n
XX6 net24 A1 ZN VPW NHVT11LL_CKT W=0.35u L=40.00n
XX2 net36 A2 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX0 A1N A1 VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX5 net24 net36 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX8 net24 A1N ZN VNW PHVT11LL_CKT W=0.35u L=40.00n
XX9 net36 A1 ZN VNW PHVT11LL_CKT W=0.35u L=40.00n
XX3 A1N A1 VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX1 net36 A2 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX4 net24 net36 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
.ENDS XNOR2V1_12TH40
.SUBCKT XNOR2V2_12TH40 A1 A2 ZN VDD VSS
XX7 net36 A1N ZN VPW NHVT11LL_CKT W=500.00n L=40.00n
XX6 net24 A1 ZN VPW NHVT11LL_CKT W=500.00n L=40.00n
XX2 net36 A2 VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX0 A1N A1 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX5 net24 net36 VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX8 net24 A1N ZN VNW PHVT11LL_CKT W=500.00n L=40.00n
XX9 net36 A1 ZN VNW PHVT11LL_CKT W=500.00n L=40.00n
XX3 A1N A1 VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX1 net36 A2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX4 net24 net36 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS XNOR2V2_12TH40
.SUBCKT XNOR2V3_12TH40 A1 A2 ZN VDD VSS
XX7 net36 A1N ZN VPW NHVT11LL_CKT W=0.7u L=40.00n
XX6 net24 A1 ZN VPW NHVT11LL_CKT W=0.7u L=40.00n
XX2 net36 A2 VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX0 A1N A1 VSS VPW NHVT11LL_CKT W=0.48u L=40.00n
XX5 net24 net36 VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX8 net24 A1N ZN VNW PHVT11LL_CKT W=0.7u L=40.00n
XX9 net36 A1 ZN VNW PHVT11LL_CKT W=0.7u L=40.00n
XX3 A1N A1 VDD VNW PHVT11LL_CKT W=0.55u L=40.00n
XX1 net36 A2 VDD VNW PHVT11LL_CKT W=0.7u L=40.00n
XX4 net24 net36 VDD VNW PHVT11LL_CKT W=0.7u L=40.00n
.ENDS XNOR2V3_12TH40
.SUBCKT XNOR2V4_12TH40 A1 A2 ZN VDD VSS
XX7 net36 A1N ZN VPW NHVT11LL_CKT W=1u L=40.00n
XX6 net24 A1 ZN VPW NHVT11LL_CKT W=1u L=40.00n
XX2 net36 A2 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX0 A1N A1 VSS VPW NHVT11LL_CKT W=0.62u L=40.00n
XX5 net24 net36 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX8 net24 A1N ZN VNW PHVT11LL_CKT W=1u L=40.00n
XX9 net36 A1 ZN VNW PHVT11LL_CKT W=1u L=40.00n
XX3 A1N A1 VDD VNW PHVT11LL_CKT W=0.71u L=40.00n
XX1 net36 A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX4 net24 net36 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS XNOR2V4_12TH40
.SUBCKT XNOR2V6_12TH40 A1 A2 ZN VDD VSS
XX7 net36 A1N ZN VPW NHVT11LL_CKT W=1.5u L=40.00n
XX6 net24 A1 ZN VPW NHVT11LL_CKT W=1.5u L=40.00n
XX2 net36 A2 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX0 A1N A1 VSS VPW NHVT11LL_CKT W=0.88u L=40.00n
XX5 net24 net36 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX8 net24 A1N ZN VNW PHVT11LL_CKT W=1.5u L=40.00n
XX9 net36 A1 ZN VNW PHVT11LL_CKT W=1.5u L=40.00n
XX3 A1N A1 VDD VNW PHVT11LL_CKT W=1u L=40.00n
XX1 net36 A2 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX4 net24 net36 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS XNOR2V6_12TH40
.SUBCKT XNOR2V8_12TH40 A1 A2 ZN VDD VSS
XX7 net36 A1N ZN VPW NHVT11LL_CKT W=2u L=40.00n
XX6 net24 A1 ZN VPW NHVT11LL_CKT W=2u L=40.00n
XX2 net36 A2 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX0 A1N A1 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX5 net24 net36 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX8 net24 A1N ZN VNW PHVT11LL_CKT W=2u L=40.00n
XX9 net36 A1 ZN VNW PHVT11LL_CKT W=2u L=40.00n
XX3 A1N A1 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 net36 A2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX4 net24 net36 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS XNOR2V8_12TH40
.SUBCKT XNOR3V0_12TH40 A1 A2 A3 ZN VDD VSS
XX19 ZN net074 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX17 A3N A3 VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX12 net12 A3 net074 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX11 net12 net31 VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX13 net31 A3N net074 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX5 net16 net24 VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX0 A2N A2 VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX2 net24 A1 VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX6 net16 A2N net31 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX7 net24 A2 net31 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX20 ZN net074 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX18 A3N A3 VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX14 net12 net31 VDD VNW PHVT11LL_CKT W=0.16u L=40.00n
XX16 net12 A3N net074 VNW PHVT11LL_CKT W=0.16u L=40.00n
XX15 net31 A3 net074 VNW PHVT11LL_CKT W=0.16u L=40.00n
XX4 net16 net24 VDD VNW PHVT11LL_CKT W=0.16u L=40.00n
XX1 net24 A1 VDD VNW PHVT11LL_CKT W=0.16u L=40.00n
XX3 A2N A2 VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX9 net24 A2N net31 VNW PHVT11LL_CKT W=0.16u L=40.00n
XX8 net16 A2 net31 VNW PHVT11LL_CKT W=0.16u L=40.00n
.ENDS XNOR3V0_12TH40
.SUBCKT XNOR3V1_12TH40 A1 A2 A3 ZN VDD VSS
XX19 ZN net074 VSS VPW NHVT11LL_CKT W=0.375u L=40.00n
XX17 A3N A3 VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX12 net12 A3 net074 VPW NHVT11LL_CKT W=0.16u L=40.00n
XX11 net12 net31 VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX13 net31 A3N net074 VPW NHVT11LL_CKT W=0.16u L=40.00n
XX5 net16 net24 VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX0 A2N A2 VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX2 net24 A1 VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX6 net16 A2N net31 VPW NHVT11LL_CKT W=0.16u L=40.00n
XX7 net24 A2 net31 VPW NHVT11LL_CKT W=0.16u L=40.00n
XX20 ZN net074 VDD VNW PHVT11LL_CKT W=0.47u L=40.00n
XX18 A3N A3 VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX14 net12 net31 VDD VNW PHVT11LL_CKT W=0.205u L=40.00n
XX16 net12 A3N net074 VNW PHVT11LL_CKT W=0.205u L=40.00n
XX15 net31 A3 net074 VNW PHVT11LL_CKT W=0.205u L=40.00n
XX4 net16 net24 VDD VNW PHVT11LL_CKT W=0.205u L=40.00n
XX1 net24 A1 VDD VNW PHVT11LL_CKT W=0.205u L=40.00n
XX3 A2N A2 VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX9 net24 A2N net31 VNW PHVT11LL_CKT W=0.205u L=40.00n
XX8 net16 A2 net31 VNW PHVT11LL_CKT W=0.205u L=40.00n
.ENDS XNOR3V1_12TH40
.SUBCKT XNOR3V2_12TH40 A1 A2 A3 ZN VDD VSS
XX19 ZN net074 VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX17 A3N A3 VSS VPW NHVT11LL_CKT W=0.345u L=40.00n
XX12 net12 A3 net074 VPW NHVT11LL_CKT W=220.00n L=40.00n
XX11 net12 net31 VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX13 net31 A3N net074 VPW NHVT11LL_CKT W=220.00n L=40.00n
XX5 net16 net24 VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX0 A2N A2 VSS VPW NHVT11LL_CKT W=340.00n L=40.00n
XX2 net24 A1 VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX6 net16 A2N net31 VPW NHVT11LL_CKT W=220.00n L=40.00n
XX7 net24 A2 net31 VPW NHVT11LL_CKT W=220.00n L=40.00n
XX20 ZN net074 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX18 A3N A3 VDD VNW PHVT11LL_CKT W=385.00n L=40.00n
XX14 net12 net31 VDD VNW PHVT11LL_CKT W=280.00n L=40.00n
XX16 net12 A3N net074 VNW PHVT11LL_CKT W=280.00n L=40.00n
XX15 net31 A3 net074 VNW PHVT11LL_CKT W=280.00n L=40.00n
XX4 net16 net24 VDD VNW PHVT11LL_CKT W=280.00n L=40.00n
XX1 net24 A1 VDD VNW PHVT11LL_CKT W=280.00n L=40.00n
XX3 A2N A2 VDD VNW PHVT11LL_CKT W=385.00n L=40.00n
XX9 net24 A2N net31 VNW PHVT11LL_CKT W=280.00n L=40.00n
XX8 net16 A2 net31 VNW PHVT11LL_CKT W=280.00n L=40.00n
.ENDS XNOR3V2_12TH40
.SUBCKT XNOR3V3_12TH40 A1 A2 A3 ZN VDD VSS
XX19 ZN net074 VSS VPW NHVT11LL_CKT W=0.76u L=40.00n
XX17 A3N A3 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX12 net12 A3 net074 VPW NHVT11LL_CKT W=0.31u L=40.00n
XX11 net12 net31 VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX13 net31 A3N net074 VPW NHVT11LL_CKT W=0.31u L=40.00n
XX5 net16 net24 VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX0 A2N A2 VSS VPW NHVT11LL_CKT W=0.385u L=40.00n
XX2 net24 A1 VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX6 net16 A2N net31 VPW NHVT11LL_CKT W=0.31u L=40.00n
XX7 net24 A2 net31 VPW NHVT11LL_CKT W=0.31u L=40.00n
XX20 ZN net074 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX18 A3N A3 VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX14 net12 net31 VDD VNW PHVT11LL_CKT W=0.39u L=40.00n
XX16 net12 A3N net074 VNW PHVT11LL_CKT W=0.39u L=40.00n
XX15 net31 A3 net074 VNW PHVT11LL_CKT W=0.39u L=40.00n
XX4 net16 net24 VDD VNW PHVT11LL_CKT W=0.39u L=40.00n
XX1 net24 A1 VDD VNW PHVT11LL_CKT W=0.39u L=40.00n
XX3 A2N A2 VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX9 net24 A2N net31 VNW PHVT11LL_CKT W=0.39u L=40.00n
XX8 net16 A2 net31 VNW PHVT11LL_CKT W=0.39u L=40.00n
.ENDS XNOR3V3_12TH40
.SUBCKT XNOR3V4_12TH40 A1 A2 A3 ZN VDD VSS
XX19 ZN net074 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX17 A3N A3 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX12 net12 A3 net074 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX11 net12 net31 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX13 net31 A3N net074 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX5 net16 net24 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX0 A2N A2 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX2 net24 A1 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX6 net16 A2N net31 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX7 net24 A2 net31 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX20 ZN net074 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX18 A3N A3 VDD VNW PHVT11LL_CKT W=0.49u L=40.00n
XX14 net12 net31 VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX16 net12 A3N net074 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX15 net31 A3 net074 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX4 net16 net24 VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX1 net24 A1 VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX3 A2N A2 VDD VNW PHVT11LL_CKT W=0.49u L=40.00n
XX9 net24 A2N net31 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX8 net16 A2 net31 VNW PHVT11LL_CKT W=0.5u L=40.00n
.ENDS XNOR3V4_12TH40
.SUBCKT XNOR3V6_12TH40 A1 A2 A3 ZN VDD VSS
XX19 ZN net074 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX17 A3N A3 VSS VPW NHVT11LL_CKT W=0.84u L=40.00n
XX12 net12 A3 net074 VPW NHVT11LL_CKT W=0.8u L=40.00n
XX11 net12 net31 VSS VPW NHVT11LL_CKT W=0.8u L=40.00n
XX13 net31 A3N net074 VPW NHVT11LL_CKT W=0.8u L=40.00n
XX5 net16 net24 VSS VPW NHVT11LL_CKT W=0.8u L=40.00n
XX0 A2N A2 VSS VPW NHVT11LL_CKT W=0.84u L=40.00n
XX2 net24 A1 VSS VPW NHVT11LL_CKT W=0.8u L=40.00n
XX6 net16 A2N net31 VPW NHVT11LL_CKT W=0.8u L=40.00n
XX7 net24 A2 net31 VPW NHVT11LL_CKT W=0.8u L=40.00n
XX20 ZN net074 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX18 A3N A3 VDD VNW PHVT11LL_CKT W=0.95u L=40.00n
XX14 net12 net31 VDD VNW PHVT11LL_CKT W=1u L=40.00n
XX16 net12 A3N net074 VNW PHVT11LL_CKT W=1u L=40.00n
XX15 net31 A3 net074 VNW PHVT11LL_CKT W=1u L=40.00n
XX4 net16 net24 VDD VNW PHVT11LL_CKT W=1u L=40.00n
XX1 net24 A1 VDD VNW PHVT11LL_CKT W=1u L=40.00n
XX3 A2N A2 VDD VNW PHVT11LL_CKT W=0.95u L=40.00n
XX9 net24 A2N net31 VNW PHVT11LL_CKT W=1u L=40.00n
XX8 net16 A2 net31 VNW PHVT11LL_CKT W=1u L=40.00n
.ENDS XNOR3V6_12TH40
.SUBCKT XNOR3V8_12TH40 A1 A2 A3 ZN VDD VSS
XX19 ZN net074 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX17 A3N A3 VSS VPW NHVT11LL_CKT W=1.04u L=40.00n
XX12 net12 A3 net074 VPW NHVT11LL_CKT W=1.2u L=40.00n
XX11 net12 net31 VSS VPW NHVT11LL_CKT W=1.2u L=40.00n
XX13 net31 A3N net074 VPW NHVT11LL_CKT W=1.2u L=40.00n
XX5 net16 net24 VSS VPW NHVT11LL_CKT W=1.2u L=40.00n
XX0 A2N A2 VSS VPW NHVT11LL_CKT W=1.04u L=40.00n
XX2 net24 A1 VSS VPW NHVT11LL_CKT W=1.2u L=40.00n
XX6 net16 A2N net31 VPW NHVT11LL_CKT W=1.2u L=40.00n
XX7 net24 A2 net31 VPW NHVT11LL_CKT W=1.2u L=40.00n
XX20 ZN net074 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX18 A3N A3 VDD VNW PHVT11LL_CKT W=1.19u L=40.00n
XX14 net12 net31 VDD VNW PHVT11LL_CKT W=1.5u L=40.00n
XX16 net12 A3N net074 VNW PHVT11LL_CKT W=1.5u L=40.00n
XX15 net31 A3 net074 VNW PHVT11LL_CKT W=1.5u L=40.00n
XX4 net16 net24 VDD VNW PHVT11LL_CKT W=1.5u L=40.00n
XX1 net24 A1 VDD VNW PHVT11LL_CKT W=1.5u L=40.00n
XX3 A2N A2 VDD VNW PHVT11LL_CKT W=1.19u L=40.00n
XX9 net24 A2N net31 VNW PHVT11LL_CKT W=1.5u L=40.00n
XX8 net16 A2 net31 VNW PHVT11LL_CKT W=1.5u L=40.00n
.ENDS XNOR3V8_12TH40
.SUBCKT XNOR4V1_12TH40 A1 A2 A3 A4 ZN VDD VSS
XX25 a3nn a3n VSS VPW NHVT11LL_CKT W=280.00n L=40.00n
XX23 a4n A4 VSS VPW NHVT11LL_CKT W=280.00n L=40.00n
XX10 a3n A3 VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX11 a2n A2 VSS VPW NHVT11LL_CKT W=280.00n L=40.00n
XX12 a1n A1 VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX13 a1nn a1n VSS VPW NHVT11LL_CKT W=280.00n L=40.00n
XX15 ZN xa1a2a3a4 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX17 xna1a2 xa3a4 xa1a2a3a4 VPW NHVT11LL_CKT W=280.00n L=40.00n
XX16 xa1a2 xna3a4 xa1a2a3a4 VPW NHVT11LL_CKT W=280.00n L=40.00n
XX33 a3n A4 xa3a4 VPW NHVT11LL_CKT W=280.00n L=40.00n
XX32 a3nn a4n xa3a4 VPW NHVT11LL_CKT W=280.00n L=40.00n
XX31 a3n a4n xna3a4 VPW NHVT11LL_CKT W=280.00n L=40.00n
XX30 a3nn A4 xna3a4 VPW NHVT11LL_CKT W=280.00n L=40.00n
XX18 a1nn A2 xna1a2 VPW NHVT11LL_CKT W=280.00n L=40.00n
XX19 a1n a2n xna1a2 VPW NHVT11LL_CKT W=280.00n L=40.00n
XX20 a1nn a2n xa1a2 VPW NHVT11LL_CKT W=280.00n L=40.00n
XX21 a1n A2 xa1a2 VPW NHVT11LL_CKT W=280.00n L=40.00n
XX24 a3nn a3n VDD VNW PHVT11LL_CKT W=350.00n L=40.00n
XX4 a4n A4 VDD VNW PHVT11LL_CKT W=350.00n L=40.00n
XX0 a2n A2 VDD VNW PHVT11LL_CKT W=350.00n L=40.00n
XX1 a3n A3 VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
XX2 a1n A1 VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
XX3 a1nn a1n VDD VNW PHVT11LL_CKT W=350.00n L=40.00n
XX5 ZN xa1a2a3a4 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX6 xna1a2 xna3a4 xa1a2a3a4 VNW PHVT11LL_CKT W=350.00n L=40.00n
XX7 xa1a2 xa3a4 xa1a2a3a4 VNW PHVT11LL_CKT W=350.00n L=40.00n
XX29 a3n a4n xa3a4 VNW PHVT11LL_CKT W=350.00n L=40.00n
XX28 a3nn A4 xa3a4 VNW PHVT11LL_CKT W=350.00n L=40.00n
XX27 a3n A4 xna3a4 VNW PHVT11LL_CKT W=350.00n L=40.00n
XX26 a3nn a4n xna3a4 VNW PHVT11LL_CKT W=350.00n L=40.00n
XX8 a1nn a2n xna1a2 VNW PHVT11LL_CKT W=350.00n L=40.00n
XX9 a1n A2 xna1a2 VNW PHVT11LL_CKT W=350.00n L=40.00n
XX14 a1nn A2 xa1a2 VNW PHVT11LL_CKT W=350.00n L=40.00n
XX22 a1n a2n xa1a2 VNW PHVT11LL_CKT W=350.00n L=40.00n
.ENDS XNOR4V1_12TH40
.SUBCKT XNOR4V2_12TH40 A1 A2 A3 A4 ZN VDD VSS
XX25 a3nn a3n VSS VPW NHVT11LL_CKT W=340.00n L=40.00n
XX23 a4n A4 VSS VPW NHVT11LL_CKT W=340.00n L=40.00n
XX10 a3n A3 VSS VPW NHVT11LL_CKT W=480.00n L=40.00n
XX11 a2n A2 VSS VPW NHVT11LL_CKT W=340.00n L=40.00n
XX12 a1n A1 VSS VPW NHVT11LL_CKT W=480.00n L=40.00n
XX13 a1nn a1n VSS VPW NHVT11LL_CKT W=340.00n L=40.00n
XX15 ZN xa1a2a3a4 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX17 xna1a2 xa3a4 xa1a2a3a4 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX16 xa1a2 xna3a4 xa1a2a3a4 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX33 a3n A4 xa3a4 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX32 a3nn a4n xa3a4 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX31 a3n a4n xna3a4 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX30 a3nn A4 xna3a4 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX18 a1nn A2 xna1a2 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX19 a1n a2n xna1a2 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX20 a1nn a2n xa1a2 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX21 a1n A2 xa1a2 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX24 a3nn a3n VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX4 a4n A4 VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX0 a2n A2 VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX1 a3n A3 VDD VNW PHVT11LL_CKT W=600.00n L=40.00n
XX2 a1n A1 VDD VNW PHVT11LL_CKT W=600.00n L=40.00n
XX3 a1nn a1n VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX5 ZN xa1a2a3a4 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX6 xna1a2 xna3a4 xa1a2a3a4 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX7 xa1a2 xa3a4 xa1a2a3a4 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX29 a3n a4n xa3a4 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX28 a3nn A4 xa3a4 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX27 a3n A4 xna3a4 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX26 a3nn a4n xna3a4 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX8 a1nn a2n xna1a2 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX9 a1n A2 xna1a2 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX14 a1nn A2 xa1a2 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX22 a1n a2n xa1a2 VNW PHVT11LL_CKT W=420.00n L=40.00n
.ENDS XNOR4V2_12TH40
.SUBCKT XNOR4V4_12TH40 A1 A2 A3 A4 ZN VDD VSS
XX25 a3nn a3n VSS VPW NHVT11LL_CKT W=690.00n L=40.00n
XX23 a4n A4 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX10 a3n A3 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX11 a2n A2 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX12 a1n A1 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX13 a1nn a1n VSS VPW NHVT11LL_CKT W=690.00n L=40.00n
XX15 ZN xa1a2a3a4 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX17 xna1a2 xa3a4 xa1a2a3a4 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX16 xa1a2 xna3a4 xa1a2a3a4 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX33 a3n A4 xa3a4 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX32 a3nn a4n xa3a4 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX31 a3n a4n xna3a4 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX30 a3nn A4 xna3a4 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX18 a1nn A2 xna1a2 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX19 a1n a2n xna1a2 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX20 a1nn a2n xa1a2 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX21 a1n A2 xa1a2 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX24 a3nn a3n VDD VNW PHVT11LL_CKT W=870.00n L=40.00n
XX4 a4n A4 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX0 a2n A2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX1 a3n A3 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX2 a1n A1 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX3 a1nn a1n VDD VNW PHVT11LL_CKT W=870.00n L=40.00n
XX5 ZN xa1a2a3a4 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX6 xna1a2 xna3a4 xa1a2a3a4 VNW PHVT11LL_CKT W=870.00n L=40.00n
XX7 xa1a2 xa3a4 xa1a2a3a4 VNW PHVT11LL_CKT W=870.00n L=40.00n
XX29 a3n a4n xa3a4 VNW PHVT11LL_CKT W=870.00n L=40.00n
XX28 a3nn A4 xa3a4 VNW PHVT11LL_CKT W=870.00n L=40.00n
XX27 a3n A4 xna3a4 VNW PHVT11LL_CKT W=870.00n L=40.00n
XX26 a3nn a4n xna3a4 VNW PHVT11LL_CKT W=870.00n L=40.00n
XX8 a1nn a2n xna1a2 VNW PHVT11LL_CKT W=870.00n L=40.00n
XX9 a1n A2 xna1a2 VNW PHVT11LL_CKT W=870.00n L=40.00n
XX14 a1nn A2 xa1a2 VNW PHVT11LL_CKT W=870.00n L=40.00n
XX22 a1n a2n xa1a2 VNW PHVT11LL_CKT W=870.00n L=40.00n
.ENDS XNOR4V4_12TH40
.SUBCKT XNOR4V8_12TH40 A1 A2 A3 A4 ZN VDD VSS
XX25 a3nn a3n VSS VPW NHVT11LL_CKT W=970.00n L=40.00n
XX23 a4n A4 VSS VPW NHVT11LL_CKT W=970.00n L=40.00n
XX10 a3n A3 VSS VPW NHVT11LL_CKT W=1.455u L=40.00n
XX11 a2n A2 VSS VPW NHVT11LL_CKT W=970.00n L=40.00n
XX12 a1n A1 VSS VPW NHVT11LL_CKT W=1.455u L=40.00n
XX13 a1nn a1n VSS VPW NHVT11LL_CKT W=970.00n L=40.00n
XX15 ZN xa1a2a3a4 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX17 xna1a2 xa3a4 xa1a2a3a4 VPW NHVT11LL_CKT W=970.00n L=40.00n
XX16 xa1a2 xna3a4 xa1a2a3a4 VPW NHVT11LL_CKT W=970.00n L=40.00n
XX33 a3n A4 xa3a4 VPW NHVT11LL_CKT W=970.00n L=40.00n
XX32 a3nn a4n xa3a4 VPW NHVT11LL_CKT W=970.00n L=40.00n
XX31 a3n a4n xna3a4 VPW NHVT11LL_CKT W=970.00n L=40.00n
XX30 a3nn A4 xna3a4 VPW NHVT11LL_CKT W=970.00n L=40.00n
XX18 a1nn A2 xna1a2 VPW NHVT11LL_CKT W=970.00n L=40.00n
XX19 a1n a2n xna1a2 VPW NHVT11LL_CKT W=970.00n L=40.00n
XX20 a1nn a2n xa1a2 VPW NHVT11LL_CKT W=970.00n L=40.00n
XX21 a1n A2 xa1a2 VPW NHVT11LL_CKT W=970.00n L=40.00n
XX24 a3nn a3n VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX4 a4n A4 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 a2n A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 a3n A3 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX2 a1n A1 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX3 a1nn a1n VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX5 ZN xa1a2a3a4 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX6 xna1a2 xna3a4 xa1a2a3a4 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX7 xa1a2 xa3a4 xa1a2a3a4 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX29 a3n a4n xa3a4 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX28 a3nn A4 xa3a4 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX27 a3n A4 xna3a4 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX26 a3nn a4n xna3a4 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX8 a1nn a2n xna1a2 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX9 a1n A2 xna1a2 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX14 a1nn A2 xa1a2 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX22 a1n a2n xa1a2 VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS XNOR4V8_12TH40
.SUBCKT XOR2V0_12TH40 A1 A2 Z VDD VSS
XX0 A1N A1 VSS VPW NHVT11LL_CKT W=0.23u L=40.00n
XX2 net8 A2 VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX6 net20 A1N Z VPW NHVT11LL_CKT W=0.25u L=40.00n
XX7 net8 A1 Z VPW NHVT11LL_CKT W=0.25u L=40.00n
XX5 net20 net8 VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX3 A1N A1 VDD VNW PHVT11LL_CKT W=0.26u L=40.00n
XX1 net8 A2 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
XX8 net20 A1 Z VNW PHVT11LL_CKT W=0.25u L=40.00n
XX9 net8 A1N Z VNW PHVT11LL_CKT W=0.25u L=40.00n
XX4 net20 net8 VDD VNW PHVT11LL_CKT W=0.305u L=40.00n
.ENDS XOR2V0_12TH40
.SUBCKT XOR2V1_12TH40 A1 A2 Z VDD VSS
XX0 A1N A1 VSS VPW NHVT11LL_CKT W=0.28u L=40.00n
XX2 net8 A2 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX6 net20 A1N Z VPW NHVT11LL_CKT W=0.35u L=40.00n
XX7 net8 A1 Z VPW NHVT11LL_CKT W=0.35u L=40.00n
XX5 net20 net8 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX3 A1N A1 VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX1 net8 A2 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
XX8 net20 A1 Z VNW PHVT11LL_CKT W=0.35u L=40.00n
XX9 net8 A1N Z VNW PHVT11LL_CKT W=0.35u L=40.00n
XX4 net20 net8 VDD VNW PHVT11LL_CKT W=0.43u L=40.00n
.ENDS XOR2V1_12TH40
.SUBCKT XOR2V2_12TH40 A1 A2 Z VDD VSS
XX0 A1N A1 VSS VPW NHVT11LL_CKT W=350.00n L=40.00n
XX2 net8 A2 VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX6 net20 A1N Z VPW NHVT11LL_CKT W=500.00n L=40.00n
XX7 net8 A1 Z VPW NHVT11LL_CKT W=500.00n L=40.00n
XX5 net20 net8 VSS VPW NHVT11LL_CKT W=500.00n L=40.00n
XX3 A1N A1 VDD VNW PHVT11LL_CKT W=400.00n L=40.00n
XX1 net8 A2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX8 net20 A1 Z VNW PHVT11LL_CKT W=500.00n L=40.00n
XX9 net8 A1N Z VNW PHVT11LL_CKT W=500.00n L=40.00n
XX4 net20 net8 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
.ENDS XOR2V2_12TH40
.SUBCKT XOR2V3_12TH40 A1 A2 Z VDD VSS
XX0 A1N A1 VSS VPW NHVT11LL_CKT W=0.48u L=40.00n
XX2 net8 A2 VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX6 net20 A1N Z VPW NHVT11LL_CKT W=0.7u L=40.00n
XX7 net8 A1 Z VPW NHVT11LL_CKT W=0.7u L=40.00n
XX5 net20 net8 VSS VPW NHVT11LL_CKT W=0.61u L=40.00n
XX3 A1N A1 VDD VNW PHVT11LL_CKT W=0.55u L=40.00n
XX1 net8 A2 VDD VNW PHVT11LL_CKT W=0.7u L=40.00n
XX8 net20 A1 Z VNW PHVT11LL_CKT W=0.7u L=40.00n
XX9 net8 A1N Z VNW PHVT11LL_CKT W=0.7u L=40.00n
XX4 net20 net8 VDD VNW PHVT11LL_CKT W=0.7u L=40.00n
.ENDS XOR2V3_12TH40
.SUBCKT XOR2V4_12TH40 A1 A2 Z VDD VSS
XX0 A1N A1 VSS VPW NHVT11LL_CKT W=0.62u L=40.00n
XX2 net8 A2 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX6 net20 A1N Z VPW NHVT11LL_CKT W=1u L=40.00n
XX7 net8 A1 Z VPW NHVT11LL_CKT W=1u L=40.00n
XX5 net20 net8 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX3 A1N A1 VDD VNW PHVT11LL_CKT W=0.71u L=40.00n
XX1 net8 A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX8 net20 A1 Z VNW PHVT11LL_CKT W=1u L=40.00n
XX9 net8 A1N Z VNW PHVT11LL_CKT W=1u L=40.00n
XX4 net20 net8 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS XOR2V4_12TH40
.SUBCKT XOR2V6_12TH40 A1 A2 Z VDD VSS
XX0 A1N A1 VSS VPW NHVT11LL_CKT W=0.88u L=40.00n
XX2 net8 A2 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX6 net20 A1N Z VPW NHVT11LL_CKT W=1.5u L=40.00n
XX7 net8 A1 Z VPW NHVT11LL_CKT W=1.5u L=40.00n
XX5 net20 net8 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX3 A1N A1 VDD VNW PHVT11LL_CKT W=1u L=40.00n
XX1 net8 A2 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX8 net20 A1 Z VNW PHVT11LL_CKT W=1.5u L=40.00n
XX9 net8 A1N Z VNW PHVT11LL_CKT W=1.5u L=40.00n
XX4 net20 net8 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
.ENDS XOR2V6_12TH40
.SUBCKT XOR2V8_12TH40 A1 A2 Z VDD VSS
XX0 A1N A1 VSS VPW NHVT11LL_CKT W=1.07u L=40.00n
XX2 net8 A2 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX6 net20 A1N Z VPW NHVT11LL_CKT W=2u L=40.00n
XX7 net8 A1 Z VPW NHVT11LL_CKT W=2u L=40.00n
XX5 net20 net8 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX3 A1N A1 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 net8 A2 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX8 net20 A1 Z VNW PHVT11LL_CKT W=2u L=40.00n
XX9 net8 A1N Z VNW PHVT11LL_CKT W=2u L=40.00n
XX4 net20 net8 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
.ENDS XOR2V8_12TH40
.SUBCKT XOR3V0_12TH40 A1 A2 A3 Z VDD VSS
XX19 Z net76 VSS VPW NHVT11LL_CKT W=0.27u L=40.00n
XX7 net57 A2 net56 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX6 net65 A2N net56 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX2 net57 A1 VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX0 A2N A2 VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX5 net65 net57 VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX11 net69 net56 VSS VPW NHVT11LL_CKT W=0.13u L=40.00n
XX12 net69 A3N net76 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX13 net56 A3 net76 VPW NHVT11LL_CKT W=0.13u L=40.00n
XX17 A3N A3 VSS VPW NHVT11LL_CKT W=0.29u L=40.00n
XX10 Z net76 VDD VNW PHVT11LL_CKT W=0.31u L=40.00n
XX8 net65 A2 net56 VNW PHVT11LL_CKT W=0.16u L=40.00n
XX9 net57 A2N net56 VNW PHVT11LL_CKT W=0.16u L=40.00n
XX3 A2N A2 VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
XX1 net57 A1 VDD VNW PHVT11LL_CKT W=0.16u L=40.00n
XX4 net65 net57 VDD VNW PHVT11LL_CKT W=0.16u L=40.00n
XX14 net69 net56 VDD VNW PHVT11LL_CKT W=0.16u L=40.00n
XX15 net56 A3N net76 VNW PHVT11LL_CKT W=0.16u L=40.00n
XX16 net69 A3 net76 VNW PHVT11LL_CKT W=0.16u L=40.00n
XX18 A3N A3 VDD VNW PHVT11LL_CKT W=0.33u L=40.00n
.ENDS XOR3V0_12TH40
.SUBCKT XOR3V1_12TH40 A1 A2 A3 Z VDD VSS
XX19 Z net76 VSS VPW NHVT11LL_CKT W=0.38u L=40.00n
XX7 net57 A2 net56 VPW NHVT11LL_CKT W=0.16u L=40.00n
XX6 net65 A2N net56 VPW NHVT11LL_CKT W=0.16u L=40.00n
XX2 net57 A1 VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX0 A2N A2 VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX5 net65 net57 VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX11 net69 net56 VSS VPW NHVT11LL_CKT W=0.16u L=40.00n
XX12 net69 A3N net76 VPW NHVT11LL_CKT W=0.16u L=40.00n
XX13 net56 A3 net76 VPW NHVT11LL_CKT W=0.16u L=40.00n
XX17 A3N A3 VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX10 Z net76 VDD VNW PHVT11LL_CKT W=0.47u L=40.00n
XX8 net65 A2 net56 VNW PHVT11LL_CKT W=0.205u L=40.00n
XX9 net57 A2N net56 VNW PHVT11LL_CKT W=0.205u L=40.00n
XX3 A2N A2 VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
XX1 net57 A1 VDD VNW PHVT11LL_CKT W=0.205u L=40.00n
XX4 net65 net57 VDD VNW PHVT11LL_CKT W=0.205u L=40.00n
XX14 net69 net56 VDD VNW PHVT11LL_CKT W=0.205u L=40.00n
XX15 net56 A3N net76 VNW PHVT11LL_CKT W=0.205u L=40.00n
XX16 net69 A3 net76 VNW PHVT11LL_CKT W=0.205u L=40.00n
XX18 A3N A3 VDD VNW PHVT11LL_CKT W=0.35u L=40.00n
.ENDS XOR3V1_12TH40
.SUBCKT XOR3V2_12TH40 A1 A2 A3 Z VDD VSS
XX19 Z net76 VSS VPW NHVT11LL_CKT W=0.54u L=40.00n
XX7 net57 A2 net56 VPW NHVT11LL_CKT W=220.00n L=40.00n
XX6 net65 A2N net56 VPW NHVT11LL_CKT W=220.00n L=40.00n
XX2 net57 A1 VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX0 A2N A2 VSS VPW NHVT11LL_CKT W=340.00n L=40.00n
XX5 net65 net57 VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX11 net69 net56 VSS VPW NHVT11LL_CKT W=220.00n L=40.00n
XX12 net69 A3N net76 VPW NHVT11LL_CKT W=220.00n L=40.00n
XX13 net56 A3 net76 VPW NHVT11LL_CKT W=220.00n L=40.00n
XX17 A3N A3 VSS VPW NHVT11LL_CKT W=340.00n L=40.00n
XX10 Z net76 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX8 net65 A2 net56 VNW PHVT11LL_CKT W=280.00n L=40.00n
XX9 net57 A2N net56 VNW PHVT11LL_CKT W=280.00n L=40.00n
XX3 A2N A2 VDD VNW PHVT11LL_CKT W=385.00n L=40.00n
XX1 net57 A1 VDD VNW PHVT11LL_CKT W=280.00n L=40.00n
XX4 net65 net57 VDD VNW PHVT11LL_CKT W=280.00n L=40.00n
XX14 net69 net56 VDD VNW PHVT11LL_CKT W=280.00n L=40.00n
XX15 net56 A3N net76 VNW PHVT11LL_CKT W=280.00n L=40.00n
XX16 net69 A3 net76 VNW PHVT11LL_CKT W=280.00n L=40.00n
XX18 A3N A3 VDD VNW PHVT11LL_CKT W=385.00n L=40.00n
.ENDS XOR3V2_12TH40
.SUBCKT XOR3V3_12TH40 A1 A2 A3 Z VDD VSS
XX19 Z net76 VSS VPW NHVT11LL_CKT W=0.76u L=40.00n
XX7 net57 A2 net56 VPW NHVT11LL_CKT W=0.31u L=40.00n
XX6 net65 A2N net56 VPW NHVT11LL_CKT W=0.31u L=40.00n
XX2 net57 A1 VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX0 A2N A2 VSS VPW NHVT11LL_CKT W=0.385u L=40.00n
XX5 net65 net57 VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX11 net69 net56 VSS VPW NHVT11LL_CKT W=0.31u L=40.00n
XX12 net69 A3N net76 VPW NHVT11LL_CKT W=0.31u L=40.00n
XX13 net56 A3 net76 VPW NHVT11LL_CKT W=0.31u L=40.00n
XX17 A3N A3 VSS VPW NHVT11LL_CKT W=0.385u L=40.00n
XX10 Z net76 VDD VNW PHVT11LL_CKT W=0.86u L=40.00n
XX8 net65 A2 net56 VNW PHVT11LL_CKT W=0.39u L=40.00n
XX9 net57 A2N net56 VNW PHVT11LL_CKT W=0.39u L=40.00n
XX3 A2N A2 VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
XX1 net57 A1 VDD VNW PHVT11LL_CKT W=0.39u L=40.00n
XX4 net65 net57 VDD VNW PHVT11LL_CKT W=0.39u L=40.00n
XX14 net69 net56 VDD VNW PHVT11LL_CKT W=0.39u L=40.00n
XX15 net56 A3N net76 VNW PHVT11LL_CKT W=0.39u L=40.00n
XX16 net69 A3 net76 VNW PHVT11LL_CKT W=0.39u L=40.00n
XX18 A3N A3 VDD VNW PHVT11LL_CKT W=0.44u L=40.00n
.ENDS XOR3V3_12TH40
.SUBCKT XOR3V4_12TH40 A1 A2 A3 Z VDD VSS
XX19 Z net76 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX7 net57 A2 net56 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX6 net65 A2N net56 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX2 net57 A1 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX0 A2N A2 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX5 net65 net57 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX11 net69 net56 VSS VPW NHVT11LL_CKT W=0.4u L=40.00n
XX12 net69 A3N net76 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX13 net56 A3 net76 VPW NHVT11LL_CKT W=0.4u L=40.00n
XX17 A3N A3 VSS VPW NHVT11LL_CKT W=0.43u L=40.00n
XX10 Z net76 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX8 net65 A2 net56 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX9 net57 A2N net56 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX3 A2N A2 VDD VNW PHVT11LL_CKT W=0.49u L=40.00n
XX1 net57 A1 VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX4 net65 net57 VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX14 net69 net56 VDD VNW PHVT11LL_CKT W=0.5u L=40.00n
XX15 net56 A3N net76 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX16 net69 A3 net76 VNW PHVT11LL_CKT W=0.5u L=40.00n
XX18 A3N A3 VDD VNW PHVT11LL_CKT W=0.49u L=40.00n
.ENDS XOR3V4_12TH40
.SUBCKT XOR3V6_12TH40 A1 A2 A3 Z VDD VSS
XX19 Z net76 VSS VPW NHVT11LL_CKT W=1.62u L=40.00n
XX7 net57 A2 net56 VPW NHVT11LL_CKT W=0.8u L=40.00n
XX6 net65 A2N net56 VPW NHVT11LL_CKT W=0.8u L=40.00n
XX2 net57 A1 VSS VPW NHVT11LL_CKT W=0.8u L=40.00n
XX0 A2N A2 VSS VPW NHVT11LL_CKT W=0.84u L=40.00n
XX5 net65 net57 VSS VPW NHVT11LL_CKT W=0.8u L=40.00n
XX11 net69 net56 VSS VPW NHVT11LL_CKT W=0.8u L=40.00n
XX12 net69 A3N net76 VPW NHVT11LL_CKT W=0.8u L=40.00n
XX13 net56 A3 net76 VPW NHVT11LL_CKT W=0.8u L=40.00n
XX17 A3N A3 VSS VPW NHVT11LL_CKT W=0.84u L=40.00n
XX10 Z net76 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX8 net65 A2 net56 VNW PHVT11LL_CKT W=1u L=40.00n
XX9 net57 A2N net56 VNW PHVT11LL_CKT W=1u L=40.00n
XX3 A2N A2 VDD VNW PHVT11LL_CKT W=0.95u L=40.00n
XX1 net57 A1 VDD VNW PHVT11LL_CKT W=1u L=40.00n
XX4 net65 net57 VDD VNW PHVT11LL_CKT W=1u L=40.00n
XX14 net69 net56 VDD VNW PHVT11LL_CKT W=1u L=40.00n
XX15 net56 A3N net76 VNW PHVT11LL_CKT W=1u L=40.00n
XX16 net69 A3 net76 VNW PHVT11LL_CKT W=1u L=40.00n
XX18 A3N A3 VDD VNW PHVT11LL_CKT W=0.95u L=40.00n
.ENDS XOR3V6_12TH40
.SUBCKT XOR3V8_12TH40 A1 A2 A3 Z VDD VSS
XX19 Z net76 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX7 net57 A2 net56 VPW NHVT11LL_CKT W=1.2u L=40.00n
XX6 net65 A2N net56 VPW NHVT11LL_CKT W=1.2u L=40.00n
XX2 net57 A1 VSS VPW NHVT11LL_CKT W=1.2u L=40.00n
XX0 A2N A2 VSS VPW NHVT11LL_CKT W=1.04u L=40.00n
XX5 net65 net57 VSS VPW NHVT11LL_CKT W=1.2u L=40.00n
XX11 net69 net56 VSS VPW NHVT11LL_CKT W=1.2u L=40.00n
XX12 net69 A3N net76 VPW NHVT11LL_CKT W=1.2u L=40.00n
XX13 net56 A3 net76 VPW NHVT11LL_CKT W=1.2u L=40.00n
XX17 A3N A3 VSS VPW NHVT11LL_CKT W=1.04u L=40.00n
XX10 Z net76 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX8 net65 A2 net56 VNW PHVT11LL_CKT W=1.5u L=40.00n
XX9 net57 A2N net56 VNW PHVT11LL_CKT W=1.5u L=40.00n
XX3 A2N A2 VDD VNW PHVT11LL_CKT W=1.19u L=40.00n
XX1 net57 A1 VDD VNW PHVT11LL_CKT W=1.5u L=40.00n
XX4 net65 net57 VDD VNW PHVT11LL_CKT W=1.5u L=40.00n
XX14 net69 net56 VDD VNW PHVT11LL_CKT W=1.5u L=40.00n
XX15 net56 A3N net76 VNW PHVT11LL_CKT W=1.5u L=40.00n
XX16 net69 A3 net76 VNW PHVT11LL_CKT W=1.5u L=40.00n
XX18 A3N A3 VDD VNW PHVT11LL_CKT W=1.19u L=40.00n
.ENDS XOR3V8_12TH40
.SUBCKT XOR4V1_12TH40 A1 A2 A3 A4 Z VDD VSS
XX13 a1nn a1n VSS VPW NHVT11LL_CKT W=280.00n L=40.00n
XX12 a1n A1 VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX11 a2n A2 VSS VPW NHVT11LL_CKT W=280.00n L=40.00n
XX10 a3n A3 VSS VPW NHVT11LL_CKT W=400.00n L=40.00n
XX15 Z net29 VSS VPW NHVT11LL_CKT W=380.00n L=40.00n
XX16 xa1a2 xa3a4 net29 VPW NHVT11LL_CKT W=280.00n L=40.00n
XX17 xna1a2 xna3a4 net29 VPW NHVT11LL_CKT W=280.00n L=40.00n
XX21 a1n A2 xa1a2 VPW NHVT11LL_CKT W=280.00n L=40.00n
XX20 a1nn a2n xa1a2 VPW NHVT11LL_CKT W=280.00n L=40.00n
XX19 a1n a2n xna1a2 VPW NHVT11LL_CKT W=280.00n L=40.00n
XX18 a1nn A2 xna1a2 VPW NHVT11LL_CKT W=280.00n L=40.00n
XX23 a4n A4 VSS VPW NHVT11LL_CKT W=280.00n L=40.00n
XX25 a3nn a3n VSS VPW NHVT11LL_CKT W=280.00n L=40.00n
XX30 a3nn A4 xna3a4 VPW NHVT11LL_CKT W=280.00n L=40.00n
XX31 a3n a4n xna3a4 VPW NHVT11LL_CKT W=280.00n L=40.00n
XX32 a3nn a4n xa3a4 VPW NHVT11LL_CKT W=280.00n L=40.00n
XX33 a3n A4 xa3a4 VPW NHVT11LL_CKT W=280.00n L=40.00n
XX3 a1nn a1n VDD VNW PHVT11LL_CKT W=350.00n L=40.00n
XX2 a1n A1 VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
XX1 a3n A3 VDD VNW PHVT11LL_CKT W=500.00n L=40.00n
XX0 a2n A2 VDD VNW PHVT11LL_CKT W=350.00n L=40.00n
XX5 Z net29 VDD VNW PHVT11LL_CKT W=430.00n L=40.00n
XX7 xa1a2 xna3a4 net29 VNW PHVT11LL_CKT W=350.00n L=40.00n
XX6 xna1a2 xa3a4 net29 VNW PHVT11LL_CKT W=350.00n L=40.00n
XX22 a1n a2n xa1a2 VNW PHVT11LL_CKT W=350.00n L=40.00n
XX14 a1nn A2 xa1a2 VNW PHVT11LL_CKT W=350.00n L=40.00n
XX9 a1n A2 xna1a2 VNW PHVT11LL_CKT W=350.00n L=40.00n
XX8 a1nn a2n xna1a2 VNW PHVT11LL_CKT W=350.00n L=40.00n
XX4 a4n A4 VDD VNW PHVT11LL_CKT W=350.00n L=40.00n
XX24 a3nn a3n VDD VNW PHVT11LL_CKT W=350.00n L=40.00n
XX26 a3nn a4n xna3a4 VNW PHVT11LL_CKT W=350.00n L=40.00n
XX27 a3n A4 xna3a4 VNW PHVT11LL_CKT W=350.00n L=40.00n
XX28 a3nn A4 xa3a4 VNW PHVT11LL_CKT W=350.00n L=40.00n
XX29 a3n a4n xa3a4 VNW PHVT11LL_CKT W=350.00n L=40.00n
.ENDS XOR4V1_12TH40
.SUBCKT XOR4V2_12TH40 A1 A2 A3 A4 Z VDD VSS
XX13 a1nn a1n VSS VPW NHVT11LL_CKT W=340.00n L=40.00n
XX12 a1n A1 VSS VPW NHVT11LL_CKT W=480.00n L=40.00n
XX11 a2n A2 VSS VPW NHVT11LL_CKT W=340.00n L=40.00n
XX10 a3n A3 VSS VPW NHVT11LL_CKT W=480.00n L=40.00n
XX15 Z net29 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX16 xa1a2 xa3a4 net29 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX17 xna1a2 xna3a4 net29 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX21 a1n A2 xa1a2 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX20 a1nn a2n xa1a2 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX19 a1n a2n xna1a2 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX18 a1nn A2 xna1a2 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX23 a4n A4 VSS VPW NHVT11LL_CKT W=340.00n L=40.00n
XX25 a3nn a3n VSS VPW NHVT11LL_CKT W=340.00n L=40.00n
XX30 a3nn A4 xna3a4 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX31 a3n a4n xna3a4 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX32 a3nn a4n xa3a4 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX33 a3n A4 xa3a4 VPW NHVT11LL_CKT W=340.00n L=40.00n
XX3 a1nn a1n VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX2 a1n A1 VDD VNW PHVT11LL_CKT W=600.00n L=40.00n
XX1 a3n A3 VDD VNW PHVT11LL_CKT W=600.00n L=40.00n
XX0 a2n A2 VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX5 Z net29 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX7 xa1a2 xna3a4 net29 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX6 xna1a2 xa3a4 net29 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX22 a1n a2n xa1a2 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX14 a1nn A2 xa1a2 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX9 a1n A2 xna1a2 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX8 a1nn a2n xna1a2 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX4 a4n A4 VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX24 a3nn a3n VDD VNW PHVT11LL_CKT W=420.00n L=40.00n
XX26 a3nn a4n xna3a4 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX27 a3n A4 xna3a4 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX28 a3nn A4 xa3a4 VNW PHVT11LL_CKT W=420.00n L=40.00n
XX29 a3n a4n xa3a4 VNW PHVT11LL_CKT W=420.00n L=40.00n
.ENDS XOR4V2_12TH40
.SUBCKT XOR4V4_12TH40 A1 A2 A3 A4 Z VDD VSS
XX13 a1nn a1n VSS VPW NHVT11LL_CKT W=690.00n L=40.00n
XX12 a1n A1 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX11 a2n A2 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX10 a3n A3 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX15 Z net29 VSS VPW NHVT11LL_CKT W=1.08u L=40.00n
XX16 xa1a2 xa3a4 net29 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX17 xna1a2 xna3a4 net29 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX21 a1n A2 xa1a2 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX20 a1nn a2n xa1a2 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX19 a1n a2n xna1a2 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX18 a1nn A2 xna1a2 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX23 a4n A4 VSS VPW NHVT11LL_CKT W=540.00n L=40.00n
XX25 a3nn a3n VSS VPW NHVT11LL_CKT W=690.00n L=40.00n
XX30 a3nn A4 xna3a4 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX31 a3n a4n xna3a4 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX32 a3nn a4n xa3a4 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX33 a3n A4 xa3a4 VPW NHVT11LL_CKT W=690.00n L=40.00n
XX3 a1nn a1n VDD VNW PHVT11LL_CKT W=870.00n L=40.00n
XX2 a1n A1 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX1 a3n A3 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX0 a2n A2 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX5 Z net29 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX7 xa1a2 xna3a4 net29 VNW PHVT11LL_CKT W=870.00n L=40.00n
XX6 xna1a2 xa3a4 net29 VNW PHVT11LL_CKT W=870.00n L=40.00n
XX22 a1n a2n xa1a2 VNW PHVT11LL_CKT W=870.00n L=40.00n
XX14 a1nn A2 xa1a2 VNW PHVT11LL_CKT W=870.00n L=40.00n
XX9 a1n A2 xna1a2 VNW PHVT11LL_CKT W=870.00n L=40.00n
XX8 a1nn a2n xna1a2 VNW PHVT11LL_CKT W=870.00n L=40.00n
XX4 a4n A4 VDD VNW PHVT11LL_CKT W=610.00n L=40.00n
XX24 a3nn a3n VDD VNW PHVT11LL_CKT W=870.00n L=40.00n
XX26 a3nn a4n xna3a4 VNW PHVT11LL_CKT W=870.00n L=40.00n
XX27 a3n A4 xna3a4 VNW PHVT11LL_CKT W=870.00n L=40.00n
XX28 a3nn A4 xa3a4 VNW PHVT11LL_CKT W=870.00n L=40.00n
XX29 a3n a4n xa3a4 VNW PHVT11LL_CKT W=870.00n L=40.00n
.ENDS XOR4V4_12TH40
.SUBCKT XOR4V8_12TH40 A1 A2 A3 A4 Z VDD VSS
XX13 a1nn a1n VSS VPW NHVT11LL_CKT W=970.00n L=40.00n
XX12 a1n A1 VSS VPW NHVT11LL_CKT W=1.455u L=40.00n
XX11 a2n A2 VSS VPW NHVT11LL_CKT W=970.00n L=40.00n
XX10 a3n A3 VSS VPW NHVT11LL_CKT W=1.455u L=40.00n
XX15 Z net29 VSS VPW NHVT11LL_CKT W=2.16u L=40.00n
XX16 xa1a2 xa3a4 net29 VPW NHVT11LL_CKT W=970.00n L=40.00n
XX17 xna1a2 xna3a4 net29 VPW NHVT11LL_CKT W=970.00n L=40.00n
XX21 a1n A2 xa1a2 VPW NHVT11LL_CKT W=970.00n L=40.00n
XX20 a1nn a2n xa1a2 VPW NHVT11LL_CKT W=970.00n L=40.00n
XX19 a1n a2n xna1a2 VPW NHVT11LL_CKT W=970.00n L=40.00n
XX18 a1nn A2 xna1a2 VPW NHVT11LL_CKT W=970.00n L=40.00n
XX23 a4n A4 VSS VPW NHVT11LL_CKT W=970.00n L=40.00n
XX25 a3nn a3n VSS VPW NHVT11LL_CKT W=970.00n L=40.00n
XX30 a3nn A4 xna3a4 VPW NHVT11LL_CKT W=970.00n L=40.00n
XX31 a3n a4n xna3a4 VPW NHVT11LL_CKT W=970.00n L=40.00n
XX32 a3nn a4n xa3a4 VPW NHVT11LL_CKT W=970.00n L=40.00n
XX33 a3n A4 xa3a4 VPW NHVT11LL_CKT W=970.00n L=40.00n
XX3 a1nn a1n VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX2 a1n A1 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX1 a3n A3 VDD VNW PHVT11LL_CKT W=1.83u L=40.00n
XX0 a2n A2 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX5 Z net29 VDD VNW PHVT11LL_CKT W=2.44u L=40.00n
XX7 xa1a2 xna3a4 net29 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX6 xna1a2 xa3a4 net29 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX22 a1n a2n xa1a2 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX14 a1nn A2 xa1a2 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX9 a1n A2 xna1a2 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX8 a1nn a2n xna1a2 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX4 a4n A4 VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX24 a3nn a3n VDD VNW PHVT11LL_CKT W=1.22u L=40.00n
XX26 a3nn a4n xna3a4 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX27 a3n A4 xna3a4 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX28 a3nn A4 xa3a4 VNW PHVT11LL_CKT W=1.22u L=40.00n
XX29 a3n a4n xa3a4 VNW PHVT11LL_CKT W=1.22u L=40.00n
.ENDS XOR4V8_12TH40
